magic
tech scmos
timestamp 1732085805
<< nwell >>
rect 873 778 945 841
rect 989 745 1061 846
rect 855 555 922 618
rect 940 610 969 618
rect 939 555 969 610
rect 1071 568 1143 631
rect 1235 535 1327 680
rect 844 308 958 371
rect 1031 333 1098 396
rect 1116 333 1145 396
rect 1255 335 1327 398
rect 909 27 1095 141
rect 909 24 1087 27
<< ntransistor >>
rect 885 721 887 761
rect 906 721 908 761
rect 931 748 933 768
rect 1001 713 1003 733
rect 1022 713 1024 733
rect 1047 715 1049 735
rect 867 478 869 538
rect 888 478 890 538
rect 909 478 911 538
rect 955 525 957 545
rect 1083 511 1085 551
rect 1104 511 1106 551
rect 1129 538 1131 558
rect 1247 503 1249 523
rect 1268 503 1270 523
rect 1289 503 1291 523
rect 1313 505 1315 525
rect 856 211 858 291
rect 877 211 879 291
rect 898 211 900 291
rect 919 211 921 291
rect 944 278 946 298
rect 1043 256 1045 316
rect 1064 256 1066 316
rect 1085 256 1087 316
rect 1131 303 1133 323
rect 1267 278 1269 318
rect 1288 278 1290 318
rect 1313 305 1315 325
rect 872 127 892 129
rect 872 106 892 108
rect 872 85 892 87
rect 872 64 892 66
rect 879 39 899 41
<< ptransistor >>
rect 885 788 887 828
rect 906 788 908 828
rect 931 788 933 828
rect 1001 755 1003 835
rect 1022 755 1024 835
rect 1047 755 1049 795
rect 867 565 869 605
rect 888 565 890 605
rect 909 565 911 605
rect 955 565 957 605
rect 1083 578 1085 618
rect 1104 578 1106 618
rect 1129 578 1131 618
rect 1247 544 1249 664
rect 1268 544 1270 664
rect 1289 544 1291 664
rect 1313 545 1315 585
rect 856 318 858 358
rect 877 318 879 358
rect 898 318 900 358
rect 919 318 921 358
rect 944 318 946 358
rect 1043 343 1045 383
rect 1064 343 1066 383
rect 1085 343 1087 383
rect 1131 343 1133 383
rect 1267 345 1269 385
rect 1288 345 1290 385
rect 1313 345 1315 385
rect 919 127 1079 129
rect 919 106 1079 108
rect 919 85 1079 87
rect 919 64 1079 66
rect 919 39 959 41
<< ndiffusion >>
rect 884 721 885 761
rect 887 721 888 761
rect 905 721 906 761
rect 908 721 909 761
rect 930 748 931 768
rect 933 748 934 768
rect 1000 713 1001 733
rect 1003 713 1004 733
rect 1021 713 1022 733
rect 1024 713 1025 733
rect 1046 715 1047 735
rect 1049 715 1050 735
rect 866 478 867 538
rect 869 478 870 538
rect 887 478 888 538
rect 890 478 891 538
rect 908 478 909 538
rect 911 478 912 538
rect 954 525 955 545
rect 957 525 958 545
rect 1082 511 1083 551
rect 1085 511 1086 551
rect 1103 511 1104 551
rect 1106 511 1107 551
rect 1128 538 1129 558
rect 1131 538 1132 558
rect 1246 503 1247 523
rect 1249 503 1250 523
rect 1267 503 1268 523
rect 1270 503 1271 523
rect 1288 503 1289 523
rect 1291 503 1292 523
rect 1312 505 1313 525
rect 1315 505 1316 525
rect 855 211 856 291
rect 858 211 859 291
rect 876 211 877 291
rect 879 211 880 291
rect 897 211 898 291
rect 900 211 901 291
rect 918 211 919 291
rect 921 211 922 291
rect 943 278 944 298
rect 946 278 947 298
rect 1042 256 1043 316
rect 1045 256 1046 316
rect 1063 256 1064 316
rect 1066 256 1067 316
rect 1084 256 1085 316
rect 1087 256 1088 316
rect 1130 303 1131 323
rect 1133 303 1134 323
rect 1266 278 1267 318
rect 1269 278 1270 318
rect 1287 278 1288 318
rect 1290 278 1291 318
rect 1312 305 1313 325
rect 1315 305 1316 325
rect 872 129 892 130
rect 872 126 892 127
rect 872 108 892 109
rect 872 105 892 106
rect 872 87 892 88
rect 872 84 892 85
rect 872 66 892 67
rect 872 63 892 64
rect 879 41 899 42
rect 879 38 899 39
<< pdiffusion >>
rect 884 788 885 828
rect 887 788 888 828
rect 905 788 906 828
rect 908 788 909 828
rect 930 788 931 828
rect 933 788 934 828
rect 1000 755 1001 835
rect 1003 755 1004 835
rect 1021 755 1022 835
rect 1024 755 1025 835
rect 1046 755 1047 795
rect 1049 755 1050 795
rect 866 565 867 605
rect 869 565 870 605
rect 887 565 888 605
rect 890 565 891 605
rect 908 565 909 605
rect 911 565 912 605
rect 954 565 955 605
rect 957 565 958 605
rect 1082 578 1083 618
rect 1085 578 1086 618
rect 1103 578 1104 618
rect 1106 578 1107 618
rect 1128 578 1129 618
rect 1131 578 1132 618
rect 1246 544 1247 664
rect 1249 544 1250 664
rect 1267 544 1268 664
rect 1270 544 1271 664
rect 1288 544 1289 664
rect 1291 544 1292 664
rect 1312 545 1313 585
rect 1315 545 1316 585
rect 855 318 856 358
rect 858 318 859 358
rect 876 318 877 358
rect 879 318 880 358
rect 897 318 898 358
rect 900 318 901 358
rect 918 318 919 358
rect 921 318 922 358
rect 943 318 944 358
rect 946 318 947 358
rect 1042 343 1043 383
rect 1045 343 1046 383
rect 1063 343 1064 383
rect 1066 343 1067 383
rect 1084 343 1085 383
rect 1087 343 1088 383
rect 1130 343 1131 383
rect 1133 343 1134 383
rect 1266 345 1267 385
rect 1269 345 1270 385
rect 1287 345 1288 385
rect 1290 345 1291 385
rect 1312 345 1313 385
rect 1315 345 1316 385
rect 919 129 1079 130
rect 919 126 1079 127
rect 919 108 1079 109
rect 919 105 1079 106
rect 919 87 1079 88
rect 919 84 1079 85
rect 919 66 1079 67
rect 919 63 1079 64
rect 919 41 959 42
rect 919 38 959 39
<< ndcontact >>
rect 880 721 884 761
rect 888 721 905 761
rect 909 721 913 761
rect 926 748 930 768
rect 934 748 938 768
rect 996 713 1000 733
rect 1004 713 1008 733
rect 1017 713 1021 733
rect 1025 713 1029 733
rect 1042 715 1046 735
rect 1050 715 1054 735
rect 862 478 866 538
rect 870 478 874 538
rect 883 478 887 538
rect 891 478 895 538
rect 904 478 908 538
rect 912 478 916 538
rect 950 525 954 545
rect 958 525 962 545
rect 1078 511 1082 551
rect 1086 511 1103 551
rect 1107 511 1111 551
rect 1124 538 1128 558
rect 1132 538 1136 558
rect 1242 503 1246 523
rect 1250 503 1254 523
rect 1263 503 1267 523
rect 1271 503 1275 523
rect 1284 503 1288 523
rect 1292 503 1296 523
rect 1308 505 1312 525
rect 1316 505 1320 525
rect 851 211 855 291
rect 859 211 863 291
rect 872 211 876 291
rect 880 211 884 291
rect 893 211 897 291
rect 901 211 905 291
rect 914 211 918 291
rect 922 211 926 291
rect 939 278 943 298
rect 947 278 951 298
rect 1038 256 1042 316
rect 1046 256 1050 316
rect 1059 256 1063 316
rect 1067 256 1071 316
rect 1080 256 1084 316
rect 1088 256 1092 316
rect 1126 303 1130 323
rect 1134 303 1138 323
rect 1262 278 1266 318
rect 1270 278 1287 318
rect 1291 278 1295 318
rect 1308 305 1312 325
rect 1316 305 1320 325
rect 872 130 892 134
rect 872 122 892 126
rect 872 109 892 113
rect 872 101 892 105
rect 872 88 892 92
rect 872 80 892 84
rect 872 67 892 71
rect 872 59 892 63
rect 879 42 899 46
rect 879 34 899 38
<< pdcontact >>
rect 880 788 884 828
rect 888 788 905 828
rect 909 788 913 828
rect 926 788 930 828
rect 934 788 938 828
rect 996 755 1000 835
rect 1004 755 1008 835
rect 1017 755 1021 835
rect 1025 755 1029 835
rect 1042 755 1046 795
rect 1050 755 1054 795
rect 862 565 866 605
rect 870 565 887 605
rect 891 565 908 605
rect 912 565 916 605
rect 950 565 954 605
rect 958 565 962 605
rect 1078 578 1082 618
rect 1086 578 1103 618
rect 1107 578 1111 618
rect 1124 578 1128 618
rect 1132 578 1136 618
rect 1242 544 1246 664
rect 1250 544 1254 664
rect 1263 544 1267 664
rect 1271 544 1275 664
rect 1284 544 1288 664
rect 1292 544 1296 664
rect 1308 545 1312 585
rect 1316 545 1320 585
rect 851 318 855 358
rect 859 318 876 358
rect 880 318 897 358
rect 901 318 918 358
rect 922 318 926 358
rect 939 318 943 358
rect 947 318 951 358
rect 1038 343 1042 383
rect 1046 343 1063 383
rect 1067 343 1084 383
rect 1088 343 1092 383
rect 1126 343 1130 383
rect 1134 343 1138 383
rect 1262 345 1266 385
rect 1270 345 1287 385
rect 1291 345 1295 385
rect 1308 345 1312 385
rect 1316 345 1320 385
rect 919 130 1079 134
rect 919 122 1079 126
rect 919 109 1079 113
rect 919 101 1079 105
rect 919 88 1079 92
rect 919 80 1079 84
rect 919 67 1079 71
rect 919 59 1079 63
rect 919 42 959 46
rect 919 34 959 38
<< polysilicon >>
rect 885 828 887 832
rect 906 828 908 847
rect 1001 835 1003 838
rect 1022 835 1024 852
rect 931 828 933 832
rect 885 761 887 788
rect 906 761 908 788
rect 931 768 933 788
rect 1047 795 1049 799
rect 931 745 933 748
rect 1001 733 1003 755
rect 1022 733 1024 755
rect 1047 735 1049 755
rect 885 718 887 721
rect 906 718 908 721
rect 1001 710 1003 713
rect 1022 710 1024 713
rect 1047 712 1049 715
rect 1247 664 1249 672
rect 1268 664 1270 686
rect 1289 664 1291 696
rect 867 605 869 609
rect 888 605 890 624
rect 909 605 911 637
rect 1083 618 1085 622
rect 1104 618 1106 637
rect 1129 618 1131 622
rect 955 605 957 609
rect 867 538 869 565
rect 888 538 890 565
rect 909 538 911 565
rect 955 545 957 565
rect 1083 551 1085 578
rect 1104 551 1106 578
rect 1129 558 1131 578
rect 955 522 957 525
rect 1313 585 1315 589
rect 1129 535 1131 538
rect 1247 523 1249 544
rect 1268 523 1270 544
rect 1289 523 1291 544
rect 1313 525 1315 545
rect 1083 508 1085 511
rect 1104 508 1106 511
rect 1247 500 1249 503
rect 1268 500 1270 503
rect 1289 500 1291 503
rect 1313 502 1315 505
rect 867 474 869 478
rect 888 474 890 478
rect 909 474 911 478
rect 856 358 858 362
rect 877 358 879 377
rect 898 358 900 404
rect 919 358 921 415
rect 1043 383 1045 387
rect 1064 383 1066 404
rect 1085 383 1087 415
rect 1131 383 1133 387
rect 1267 385 1269 389
rect 1288 385 1290 404
rect 1313 385 1315 389
rect 944 358 946 362
rect 856 291 858 318
rect 877 291 879 318
rect 898 291 900 318
rect 919 291 921 318
rect 944 298 946 318
rect 1043 316 1045 343
rect 1064 316 1066 343
rect 1085 316 1087 343
rect 1131 323 1133 343
rect 944 275 946 278
rect 1267 318 1269 345
rect 1288 318 1290 345
rect 1313 325 1315 345
rect 1131 300 1133 303
rect 1313 302 1315 305
rect 1267 275 1269 278
rect 1288 275 1290 278
rect 1043 252 1045 256
rect 1064 252 1066 256
rect 1085 252 1087 256
rect 856 208 858 211
rect 877 208 879 211
rect 898 208 900 211
rect 919 208 921 211
rect 868 127 872 129
rect 892 127 919 129
rect 1079 127 1086 129
rect 868 106 872 108
rect 892 106 919 108
rect 1079 106 1101 108
rect 868 85 872 87
rect 892 85 919 87
rect 1079 85 1114 87
rect 868 64 872 66
rect 892 64 919 66
rect 1079 64 1125 66
rect 876 39 879 41
rect 899 39 919 41
rect 959 39 1086 41
<< polycontact >>
rect 1020 852 1026 857
rect 904 847 910 852
rect 878 768 885 774
rect 927 771 931 776
rect 994 736 1001 742
rect 1043 738 1047 743
rect 1287 696 1293 701
rect 1266 686 1272 691
rect 907 637 913 642
rect 1102 637 1108 642
rect 886 624 892 629
rect 860 545 867 551
rect 951 548 955 553
rect 1076 558 1083 564
rect 1125 561 1129 566
rect 1240 526 1247 532
rect 1309 528 1313 533
rect 917 415 923 420
rect 1083 415 1089 420
rect 896 404 902 409
rect 875 377 881 382
rect 1062 404 1068 409
rect 1286 404 1292 409
rect 1036 323 1043 329
rect 849 298 856 304
rect 940 301 944 306
rect 1127 326 1131 331
rect 1260 325 1267 331
rect 1309 328 1313 333
rect 899 129 905 136
rect 1101 104 1106 110
rect 1114 83 1119 89
rect 1125 62 1130 68
rect 902 41 907 45
<< metal1 >>
rect 876 876 1086 879
rect 876 871 1068 876
rect 1074 871 1086 876
rect 876 869 1061 871
rect 876 868 945 869
rect 788 847 835 852
rect 840 847 904 852
rect 937 841 945 868
rect 957 852 1020 857
rect 1053 846 1061 869
rect 873 833 945 841
rect 989 838 1061 846
rect 996 835 1000 838
rect 880 828 884 833
rect 909 828 913 833
rect 926 828 930 833
rect 788 768 844 774
rect 849 768 878 774
rect 893 769 898 788
rect 919 771 927 776
rect 934 775 938 788
rect 919 769 923 771
rect 893 765 923 769
rect 934 770 952 775
rect 934 768 938 770
rect 909 761 913 765
rect 1008 755 1017 835
rect 1042 795 1046 838
rect 926 731 930 748
rect 1025 743 1029 755
rect 952 736 994 742
rect 1009 738 1043 743
rect 1050 742 1054 755
rect 1009 733 1014 738
rect 1050 737 1149 742
rect 1050 735 1054 737
rect 919 728 930 731
rect 880 711 884 721
rect 919 711 925 728
rect 1008 713 1017 733
rect 870 709 931 711
rect 996 709 1000 713
rect 1025 709 1029 713
rect 1042 709 1046 715
rect 870 703 1006 709
rect 1013 703 1079 709
rect 1185 705 1353 713
rect 1360 705 1361 713
rect 1208 696 1287 701
rect 793 684 1046 690
rect 1024 659 1068 664
rect 1074 659 1195 664
rect 1024 656 1195 659
rect 857 648 1029 656
rect 815 637 844 642
rect 849 637 907 642
rect 913 637 1102 642
rect 1135 631 1143 656
rect 1208 650 1214 696
rect 796 624 823 629
rect 828 624 886 629
rect 1071 623 1143 631
rect 1159 646 1214 650
rect 1222 686 1266 691
rect 1078 618 1082 623
rect 1107 618 1111 623
rect 855 610 969 618
rect 862 605 866 610
rect 898 605 902 610
rect 950 605 954 610
rect 1124 618 1128 623
rect 840 545 860 551
rect 875 546 879 565
rect 912 546 916 565
rect 943 548 951 553
rect 958 552 962 565
rect 999 558 1046 564
rect 1053 558 1076 564
rect 1091 559 1096 578
rect 1117 561 1125 566
rect 1132 565 1136 578
rect 1159 565 1163 646
rect 1117 559 1121 561
rect 1091 555 1121 559
rect 1132 560 1163 565
rect 1132 558 1136 560
rect 943 546 947 548
rect 875 542 947 546
rect 958 547 1052 552
rect 1107 551 1111 555
rect 958 545 962 547
rect 912 538 916 542
rect 874 478 883 538
rect 895 478 904 538
rect 950 498 954 525
rect 1222 553 1228 686
rect 1319 680 1327 705
rect 1235 672 1327 680
rect 1242 664 1246 672
rect 1254 544 1263 664
rect 1275 544 1284 664
rect 1308 585 1312 672
rect 1124 521 1128 538
rect 1292 533 1296 544
rect 1212 526 1240 532
rect 1255 528 1309 533
rect 1316 532 1320 545
rect 1255 523 1260 528
rect 1292 523 1296 528
rect 1316 527 1375 532
rect 1316 525 1320 527
rect 1117 518 1128 521
rect 1078 498 1082 511
rect 1117 498 1121 518
rect 1254 503 1263 523
rect 1275 503 1284 523
rect 1242 498 1246 503
rect 1277 498 1281 503
rect 1308 498 1312 505
rect 950 493 1006 498
rect 1013 493 1187 498
rect 1197 493 1361 498
rect 862 467 866 478
rect 950 467 954 493
rect 853 459 954 467
rect 782 447 1206 452
rect 848 426 1167 434
rect 1176 431 1219 434
rect 1176 426 1353 431
rect 1205 423 1353 426
rect 1360 423 1361 431
rect 828 415 917 420
rect 923 415 1083 420
rect 784 404 896 409
rect 902 404 1062 409
rect 1068 404 1286 409
rect 1319 398 1327 423
rect 1031 388 1145 396
rect 1255 390 1327 398
rect 1038 383 1042 388
rect 1074 383 1078 388
rect 1126 383 1130 388
rect 1262 385 1266 390
rect 1291 385 1295 390
rect 840 377 875 382
rect 844 363 958 371
rect 851 358 855 363
rect 886 358 890 363
rect 922 358 926 363
rect 939 358 943 363
rect 1308 385 1312 390
rect 999 323 1036 329
rect 1051 324 1055 343
rect 1088 324 1092 343
rect 1119 326 1127 331
rect 1134 330 1138 343
rect 1119 324 1123 326
rect 1051 320 1123 324
rect 1134 325 1146 330
rect 1212 325 1260 331
rect 1275 326 1280 345
rect 1301 328 1309 333
rect 1316 332 1320 345
rect 1301 326 1305 328
rect 1134 323 1138 325
rect 815 298 849 304
rect 864 299 868 318
rect 907 299 911 318
rect 932 301 940 306
rect 947 305 951 318
rect 1088 316 1092 320
rect 932 299 936 301
rect 864 295 936 299
rect 947 300 983 305
rect 947 298 951 300
rect 922 291 926 295
rect 863 211 872 291
rect 884 211 893 291
rect 905 211 914 291
rect 939 223 943 278
rect 1050 256 1059 316
rect 1071 256 1080 316
rect 1275 322 1305 326
rect 1316 327 1351 332
rect 1316 325 1320 327
rect 1291 318 1295 322
rect 1126 268 1130 303
rect 1308 288 1312 305
rect 1301 285 1312 288
rect 1262 268 1266 278
rect 1301 268 1307 285
rect 1126 260 1188 268
rect 1197 260 1326 268
rect 1038 223 1042 256
rect 1126 223 1130 260
rect 939 215 1130 223
rect 851 198 855 211
rect 939 198 943 215
rect 793 190 943 198
rect 810 173 843 178
rect 853 134 861 190
rect 1348 178 1351 327
rect 899 136 905 178
rect 853 130 872 134
rect 853 99 861 130
rect 1087 134 1095 141
rect 1079 130 1095 134
rect 872 121 892 122
rect 872 116 900 121
rect 872 113 892 116
rect 872 99 892 101
rect 853 95 892 99
rect 853 63 861 95
rect 872 92 892 95
rect 872 77 892 80
rect 896 77 900 116
rect 919 113 1079 122
rect 919 92 1079 101
rect 872 73 900 77
rect 872 71 892 73
rect 896 63 900 73
rect 919 71 1079 80
rect 853 59 872 63
rect 896 59 919 63
rect 853 46 861 59
rect 896 53 900 59
rect 896 49 907 53
rect 853 42 879 46
rect 902 45 907 49
rect 1087 46 1095 130
rect 1101 110 1106 172
rect 1114 89 1119 172
rect 1125 172 1351 178
rect 1125 68 1130 172
rect 853 2 861 42
rect 959 42 1095 46
rect 899 34 919 38
rect 1087 35 1095 42
rect 1150 35 1158 148
rect 901 -3 906 34
rect 1087 24 1158 35
<< m2contact >>
rect 835 847 840 852
rect 1353 705 1360 713
rect 808 637 815 642
rect 823 624 828 629
rect 835 545 840 551
rect 993 558 999 564
rect 1052 547 1058 552
rect 1222 546 1228 553
rect 1206 526 1212 532
rect 1187 493 1197 498
rect 1206 447 1212 452
rect 1167 426 1176 434
rect 1353 423 1360 431
rect 823 415 828 420
rect 835 377 840 382
rect 993 323 999 329
rect 1146 325 1153 330
rect 1206 325 1212 331
rect 808 298 815 304
rect 983 300 989 305
rect 1188 260 1197 268
rect 1101 172 1106 178
rect 1114 172 1119 178
rect 1150 148 1158 154
<< metal2 >>
rect 808 304 815 637
rect 823 420 828 624
rect 835 551 840 847
rect 835 382 840 545
rect 993 329 999 558
rect 1052 506 1058 547
rect 1146 540 1228 546
rect 1146 506 1153 540
rect 1052 501 1153 506
rect 1188 498 1197 499
rect 983 178 989 300
rect 1146 200 1153 325
rect 1114 195 1153 200
rect 1114 178 1119 195
rect 983 172 1101 178
rect 1167 154 1176 426
rect 1188 268 1197 493
rect 1206 452 1212 526
rect 1206 331 1212 447
rect 1353 431 1360 705
rect 1158 148 1176 154
<< m3contact >>
rect 952 736 958 742
rect 1185 705 1195 713
rect 952 684 958 690
rect 1185 656 1195 664
rect 964 648 969 654
rect 964 613 969 618
rect 951 426 958 434
rect 951 363 958 371
rect 1103 426 1109 434
rect 837 173 843 178
rect 899 173 905 178
<< m123contact >>
rect 1068 871 1074 876
rect 952 851 957 857
rect 844 768 849 774
rect 952 770 957 775
rect 1006 703 1013 709
rect 1046 684 1053 690
rect 1068 659 1074 664
rect 844 637 849 642
rect 1046 558 1053 564
rect 1006 493 1013 498
<< metal3 >>
rect 952 775 957 851
rect 844 642 849 768
rect 952 690 958 736
rect 964 618 969 648
rect 1006 498 1013 703
rect 1046 564 1053 684
rect 1068 664 1074 871
rect 1185 664 1195 705
rect 951 371 958 426
rect 1103 388 1109 426
rect 843 173 899 178
<< labels >>
rlabel metal1 875 705 928 709 1 Gnd
rlabel metal1 875 705 928 709 1 GND
rlabel metal1 856 770 875 772 1 P1
rlabel metal1 880 848 899 850 1 G0
rlabel metal1 981 738 991 740 1 G1
rlabel metal1 996 873 1049 877 5 VDD
rlabel metal1 862 650 915 654 5 VDD
rlabel metal1 857 461 910 465 1 Gnd
rlabel metal1 857 461 910 465 1 GND
rlabel metal1 1078 658 1131 662 5 VDD
rlabel metal1 866 626 882 628 1 P2
rlabel metal1 1111 738 1139 741 1 C2
rlabel metal1 1242 707 1295 711 5 VDD
rlabel metal1 1220 528 1238 530 1 G2
rlabel metal1 1320 528 1344 531 1 C3
rlabel metal1 846 192 899 196 1 Gnd
rlabel metal1 846 192 899 196 1 GND
rlabel metal1 851 428 904 432 5 VDD
rlabel metal1 1038 428 1091 432 5 VDD
rlabel metal1 1033 217 1086 221 1 Gnd
rlabel metal1 1033 217 1086 221 1 GND
rlabel metal1 874 406 895 408 1 P3
rlabel metal1 1262 425 1315 429 5 VDD
rlabel metal1 1257 262 1310 266 1 Gnd
rlabel metal1 1257 262 1310 266 1 GND
rlabel metal1 1152 81 1156 134 7 VDD
rlabel metal1 855 86 859 139 3 Gnd
rlabel metal1 855 86 859 139 3 GND
rlabel metal1 901 148 903 163 1 G3
rlabel metal1 903 4 905 19 1 C4
rlabel metal1 1052 738 1059 740 1 C2
<< end >>
