magic
tech scmos
timestamp 1732102893
<< nwell >>
rect 2244 1366 2277 1403
rect 2283 1366 2309 1403
rect 2325 1366 2353 1403
rect 2370 1366 2398 1403
rect 2010 1208 2038 1245
rect 2055 1208 2083 1245
rect 2099 1208 2125 1245
rect 2131 1208 2164 1245
rect 2250 1162 2283 1199
rect 2289 1162 2315 1199
rect 2331 1162 2359 1199
rect 2376 1162 2404 1199
rect 2504 1195 2529 1252
rect 2541 1167 2566 1207
rect 2574 1200 2599 1240
rect 2617 1194 2642 1251
rect 2688 1193 2759 1256
rect 2827 1158 2852 1215
rect 2864 1130 2889 1170
rect 2897 1163 2922 1203
rect 2940 1157 2965 1214
rect 3066 1190 3091 1247
rect 3103 1162 3128 1202
rect 3136 1195 3161 1235
rect 3179 1189 3204 1246
rect 3353 1174 3386 1211
rect 3392 1174 3418 1211
rect 3434 1174 3462 1211
rect 3479 1174 3507 1211
rect 2253 1033 2286 1070
rect 2292 1033 2318 1070
rect 2334 1033 2362 1070
rect 2379 1033 2407 1070
rect 3356 1038 3389 1075
rect 3395 1038 3421 1075
rect 3437 1038 3465 1075
rect 3482 1038 3510 1075
rect 2263 872 2296 909
rect 2302 872 2328 909
rect 2344 872 2372 909
rect 2389 872 2417 909
rect 2484 901 2509 958
rect 2521 873 2546 913
rect 2554 906 2579 946
rect 2597 900 2622 957
rect 2668 899 2739 962
rect 2903 933 2975 996
rect 3019 900 3091 1001
rect 2263 747 2296 784
rect 2302 747 2328 784
rect 2344 747 2372 784
rect 2389 747 2417 784
rect 2494 656 2519 713
rect 2531 628 2556 668
rect 2564 661 2589 701
rect 2607 655 2632 712
rect 2678 654 2749 717
rect 2885 710 2952 773
rect 2970 765 2999 773
rect 2969 710 2999 765
rect 3101 723 3173 786
rect 3265 690 3357 835
rect 2263 581 2296 618
rect 2302 581 2328 618
rect 2344 581 2372 618
rect 2389 581 2417 618
rect 2263 456 2296 493
rect 2302 456 2328 493
rect 2344 456 2372 493
rect 2389 456 2417 493
rect 2874 463 2988 526
rect 3061 488 3128 551
rect 3146 488 3175 551
rect 3285 490 3357 553
rect 2509 402 2534 459
rect 2546 374 2571 414
rect 2579 407 2604 447
rect 2622 401 2647 458
rect 2693 400 2764 463
rect 2311 313 2344 350
rect 2350 313 2376 350
rect 2392 313 2420 350
rect 2437 313 2465 350
rect 2939 182 3125 296
rect 3249 217 3274 274
rect 3286 189 3311 229
rect 3319 222 3344 262
rect 3362 216 3387 273
rect 2939 179 3117 182
rect 3499 145 3532 182
rect 3538 145 3564 182
rect 3580 145 3608 182
rect 3625 145 3653 182
rect 2953 51 2986 88
rect 2992 51 3018 88
rect 3034 51 3062 88
rect 3079 51 3107 88
<< ntransistor >>
rect 2252 1340 2254 1350
rect 2288 1340 2290 1350
rect 2296 1340 2298 1350
rect 2332 1340 2334 1350
rect 2340 1340 2342 1350
rect 2383 1340 2385 1350
rect 2023 1261 2025 1271
rect 2066 1261 2068 1271
rect 2074 1261 2076 1271
rect 2110 1261 2112 1271
rect 2118 1261 2120 1271
rect 2154 1261 2156 1271
rect 2552 1217 2554 1237
rect 2515 1165 2517 1185
rect 2585 1170 2587 1190
rect 2628 1164 2630 1184
rect 2258 1136 2260 1146
rect 2294 1136 2296 1146
rect 2302 1136 2304 1146
rect 2338 1136 2340 1146
rect 2346 1136 2348 1146
rect 2389 1136 2391 1146
rect 2699 1136 2701 1176
rect 2720 1136 2722 1176
rect 2745 1163 2747 1183
rect 2875 1180 2877 1200
rect 3114 1212 3116 1232
rect 2838 1128 2840 1148
rect 2908 1133 2910 1153
rect 3077 1160 3079 1180
rect 3147 1165 3149 1185
rect 3190 1159 3192 1179
rect 3361 1148 3363 1158
rect 3397 1148 3399 1158
rect 3405 1148 3407 1158
rect 3441 1148 3443 1158
rect 3449 1148 3451 1158
rect 3492 1148 3494 1158
rect 2951 1127 2953 1147
rect 2261 1007 2263 1017
rect 2297 1007 2299 1017
rect 2305 1007 2307 1017
rect 2341 1007 2343 1017
rect 2349 1007 2351 1017
rect 2392 1007 2394 1017
rect 3364 1012 3366 1022
rect 3400 1012 3402 1022
rect 3408 1012 3410 1022
rect 3444 1012 3446 1022
rect 3452 1012 3454 1022
rect 3495 1012 3497 1022
rect 2532 923 2534 943
rect 2495 871 2497 891
rect 2565 876 2567 896
rect 2608 870 2610 890
rect 2271 846 2273 856
rect 2307 846 2309 856
rect 2315 846 2317 856
rect 2351 846 2353 856
rect 2359 846 2361 856
rect 2402 846 2404 856
rect 2679 842 2681 882
rect 2700 842 2702 882
rect 2725 869 2727 889
rect 2915 876 2917 916
rect 2936 876 2938 916
rect 2961 903 2963 923
rect 3031 868 3033 888
rect 3052 868 3054 888
rect 3077 870 3079 890
rect 2271 721 2273 731
rect 2307 721 2309 731
rect 2315 721 2317 731
rect 2351 721 2353 731
rect 2359 721 2361 731
rect 2402 721 2404 731
rect 2542 678 2544 698
rect 2505 626 2507 646
rect 2575 631 2577 651
rect 2618 625 2620 645
rect 2689 597 2691 637
rect 2710 597 2712 637
rect 2735 624 2737 644
rect 2897 633 2899 693
rect 2918 633 2920 693
rect 2939 633 2941 693
rect 2985 680 2987 700
rect 3113 666 3115 706
rect 3134 666 3136 706
rect 3159 693 3161 713
rect 3277 658 3279 678
rect 3298 658 3300 678
rect 3319 658 3321 678
rect 3343 660 3345 680
rect 2271 555 2273 565
rect 2307 555 2309 565
rect 2315 555 2317 565
rect 2351 555 2353 565
rect 2359 555 2361 565
rect 2402 555 2404 565
rect 2271 430 2273 440
rect 2307 430 2309 440
rect 2315 430 2317 440
rect 2351 430 2353 440
rect 2359 430 2361 440
rect 2402 430 2404 440
rect 2557 424 2559 444
rect 2520 372 2522 392
rect 2590 377 2592 397
rect 2633 371 2635 391
rect 2704 343 2706 383
rect 2725 343 2727 383
rect 2750 370 2752 390
rect 2886 366 2888 446
rect 2907 366 2909 446
rect 2928 366 2930 446
rect 2949 366 2951 446
rect 2974 433 2976 453
rect 3073 411 3075 471
rect 3094 411 3096 471
rect 3115 411 3117 471
rect 3161 458 3163 478
rect 3297 433 3299 473
rect 3318 433 3320 473
rect 3343 460 3345 480
rect 2319 287 2321 297
rect 2355 287 2357 297
rect 2363 287 2365 297
rect 2399 287 2401 297
rect 2407 287 2409 297
rect 2450 287 2452 297
rect 2902 282 2922 284
rect 2902 261 2922 263
rect 2902 240 2922 242
rect 3297 239 3299 259
rect 2902 219 2922 221
rect 2909 194 2929 196
rect 3260 187 3262 207
rect 3330 192 3332 212
rect 3373 186 3375 206
rect 3507 119 3509 129
rect 3543 119 3545 129
rect 3551 119 3553 129
rect 3587 119 3589 129
rect 3595 119 3597 129
rect 3638 119 3640 129
rect 2961 25 2963 35
rect 2997 25 2999 35
rect 3005 25 3007 35
rect 3041 25 3043 35
rect 3049 25 3051 35
rect 3092 25 3094 35
<< ptransistor >>
rect 2256 1372 2258 1397
rect 2264 1372 2266 1397
rect 2294 1372 2296 1397
rect 2338 1372 2340 1397
rect 2383 1372 2385 1397
rect 2023 1214 2025 1239
rect 2068 1214 2070 1239
rect 2112 1214 2114 1239
rect 2142 1214 2144 1239
rect 2150 1214 2152 1239
rect 2515 1205 2517 1245
rect 2585 1210 2587 1230
rect 2262 1168 2264 1193
rect 2270 1168 2272 1193
rect 2300 1168 2302 1193
rect 2344 1168 2346 1193
rect 2389 1168 2391 1193
rect 2628 1204 2630 1244
rect 2552 1177 2554 1197
rect 2699 1203 2701 1243
rect 2720 1203 2722 1243
rect 2745 1203 2747 1243
rect 2838 1168 2840 1208
rect 2908 1173 2910 1193
rect 2951 1167 2953 1207
rect 3077 1200 3079 1240
rect 3147 1205 3149 1225
rect 3190 1199 3192 1239
rect 2875 1140 2877 1160
rect 3114 1172 3116 1192
rect 3365 1180 3367 1205
rect 3373 1180 3375 1205
rect 3403 1180 3405 1205
rect 3447 1180 3449 1205
rect 3492 1180 3494 1205
rect 2265 1039 2267 1064
rect 2273 1039 2275 1064
rect 2303 1039 2305 1064
rect 2347 1039 2349 1064
rect 2392 1039 2394 1064
rect 3368 1044 3370 1069
rect 3376 1044 3378 1069
rect 3406 1044 3408 1069
rect 3450 1044 3452 1069
rect 3495 1044 3497 1069
rect 2495 911 2497 951
rect 2565 916 2567 936
rect 2275 878 2277 903
rect 2283 878 2285 903
rect 2313 878 2315 903
rect 2357 878 2359 903
rect 2402 878 2404 903
rect 2608 910 2610 950
rect 2532 883 2534 903
rect 2679 909 2681 949
rect 2700 909 2702 949
rect 2725 909 2727 949
rect 2915 943 2917 983
rect 2936 943 2938 983
rect 2961 943 2963 983
rect 3031 910 3033 990
rect 3052 910 3054 990
rect 3077 910 3079 950
rect 2275 753 2277 778
rect 2283 753 2285 778
rect 2313 753 2315 778
rect 2357 753 2359 778
rect 2402 753 2404 778
rect 2505 666 2507 706
rect 2575 671 2577 691
rect 2618 665 2620 705
rect 2897 720 2899 760
rect 2918 720 2920 760
rect 2939 720 2941 760
rect 2985 720 2987 760
rect 3113 733 3115 773
rect 3134 733 3136 773
rect 3159 733 3161 773
rect 2542 638 2544 658
rect 2689 664 2691 704
rect 2710 664 2712 704
rect 2735 664 2737 704
rect 2275 587 2277 612
rect 2283 587 2285 612
rect 2313 587 2315 612
rect 2357 587 2359 612
rect 2402 587 2404 612
rect 3277 699 3279 819
rect 3298 699 3300 819
rect 3319 699 3321 819
rect 3343 700 3345 740
rect 2275 462 2277 487
rect 2283 462 2285 487
rect 2313 462 2315 487
rect 2357 462 2359 487
rect 2402 462 2404 487
rect 2886 473 2888 513
rect 2907 473 2909 513
rect 2928 473 2930 513
rect 2949 473 2951 513
rect 2974 473 2976 513
rect 3073 498 3075 538
rect 3094 498 3096 538
rect 3115 498 3117 538
rect 3161 498 3163 538
rect 3297 500 3299 540
rect 3318 500 3320 540
rect 3343 500 3345 540
rect 2520 412 2522 452
rect 2590 417 2592 437
rect 2633 411 2635 451
rect 2557 384 2559 404
rect 2704 410 2706 450
rect 2725 410 2727 450
rect 2750 410 2752 450
rect 2323 319 2325 344
rect 2331 319 2333 344
rect 2361 319 2363 344
rect 2405 319 2407 344
rect 2450 319 2452 344
rect 2949 282 3109 284
rect 2949 261 3109 263
rect 2949 240 3109 242
rect 3260 227 3262 267
rect 3330 232 3332 252
rect 2949 219 3109 221
rect 3373 226 3375 266
rect 2949 194 2989 196
rect 3297 199 3299 219
rect 3511 151 3513 176
rect 3519 151 3521 176
rect 3549 151 3551 176
rect 3593 151 3595 176
rect 3638 151 3640 176
rect 2965 57 2967 82
rect 2973 57 2975 82
rect 3003 57 3005 82
rect 3047 57 3049 82
rect 3092 57 3094 82
<< ndiffusion >>
rect 2251 1340 2252 1350
rect 2254 1340 2255 1350
rect 2287 1340 2288 1350
rect 2290 1340 2291 1350
rect 2295 1340 2296 1350
rect 2298 1340 2299 1350
rect 2331 1340 2332 1350
rect 2334 1340 2335 1350
rect 2339 1340 2340 1350
rect 2342 1340 2343 1350
rect 2382 1340 2383 1350
rect 2385 1340 2386 1350
rect 2022 1261 2023 1271
rect 2025 1261 2026 1271
rect 2065 1261 2066 1271
rect 2068 1261 2069 1271
rect 2073 1261 2074 1271
rect 2076 1261 2077 1271
rect 2109 1261 2110 1271
rect 2112 1261 2113 1271
rect 2117 1261 2118 1271
rect 2120 1261 2121 1271
rect 2153 1261 2154 1271
rect 2156 1261 2157 1271
rect 2551 1217 2552 1237
rect 2554 1217 2555 1237
rect 2514 1165 2515 1185
rect 2517 1165 2518 1185
rect 2584 1170 2585 1190
rect 2587 1170 2588 1190
rect 2627 1164 2628 1184
rect 2630 1164 2631 1184
rect 2257 1136 2258 1146
rect 2260 1136 2261 1146
rect 2293 1136 2294 1146
rect 2296 1136 2297 1146
rect 2301 1136 2302 1146
rect 2304 1136 2305 1146
rect 2337 1136 2338 1146
rect 2340 1136 2341 1146
rect 2345 1136 2346 1146
rect 2348 1136 2349 1146
rect 2388 1136 2389 1146
rect 2391 1136 2392 1146
rect 2698 1136 2699 1176
rect 2701 1136 2702 1176
rect 2719 1136 2720 1176
rect 2722 1136 2723 1176
rect 2744 1163 2745 1183
rect 2747 1163 2748 1183
rect 2874 1180 2875 1200
rect 2877 1180 2878 1200
rect 3113 1212 3114 1232
rect 3116 1212 3117 1232
rect 2837 1128 2838 1148
rect 2840 1128 2841 1148
rect 2907 1133 2908 1153
rect 2910 1133 2911 1153
rect 3076 1160 3077 1180
rect 3079 1160 3080 1180
rect 3146 1165 3147 1185
rect 3149 1165 3150 1185
rect 3189 1159 3190 1179
rect 3192 1159 3193 1179
rect 3360 1148 3361 1158
rect 3363 1148 3364 1158
rect 3396 1148 3397 1158
rect 3399 1148 3400 1158
rect 3404 1148 3405 1158
rect 3407 1148 3408 1158
rect 3440 1148 3441 1158
rect 3443 1148 3444 1158
rect 3448 1148 3449 1158
rect 3451 1148 3452 1158
rect 3491 1148 3492 1158
rect 3494 1148 3495 1158
rect 2950 1127 2951 1147
rect 2953 1127 2954 1147
rect 2260 1007 2261 1017
rect 2263 1007 2264 1017
rect 2296 1007 2297 1017
rect 2299 1007 2300 1017
rect 2304 1007 2305 1017
rect 2307 1007 2308 1017
rect 2340 1007 2341 1017
rect 2343 1007 2344 1017
rect 2348 1007 2349 1017
rect 2351 1007 2352 1017
rect 2391 1007 2392 1017
rect 2394 1007 2395 1017
rect 3363 1012 3364 1022
rect 3366 1012 3367 1022
rect 3399 1012 3400 1022
rect 3402 1012 3403 1022
rect 3407 1012 3408 1022
rect 3410 1012 3411 1022
rect 3443 1012 3444 1022
rect 3446 1012 3447 1022
rect 3451 1012 3452 1022
rect 3454 1012 3455 1022
rect 3494 1012 3495 1022
rect 3497 1012 3498 1022
rect 2531 923 2532 943
rect 2534 923 2535 943
rect 2494 871 2495 891
rect 2497 871 2498 891
rect 2564 876 2565 896
rect 2567 876 2568 896
rect 2607 870 2608 890
rect 2610 870 2611 890
rect 2270 846 2271 856
rect 2273 846 2274 856
rect 2306 846 2307 856
rect 2309 846 2310 856
rect 2314 846 2315 856
rect 2317 846 2318 856
rect 2350 846 2351 856
rect 2353 846 2354 856
rect 2358 846 2359 856
rect 2361 846 2362 856
rect 2401 846 2402 856
rect 2404 846 2405 856
rect 2678 842 2679 882
rect 2681 842 2682 882
rect 2699 842 2700 882
rect 2702 842 2703 882
rect 2724 869 2725 889
rect 2727 869 2728 889
rect 2914 876 2915 916
rect 2917 876 2918 916
rect 2935 876 2936 916
rect 2938 876 2939 916
rect 2960 903 2961 923
rect 2963 903 2964 923
rect 3030 868 3031 888
rect 3033 868 3034 888
rect 3051 868 3052 888
rect 3054 868 3055 888
rect 3076 870 3077 890
rect 3079 870 3080 890
rect 2270 721 2271 731
rect 2273 721 2274 731
rect 2306 721 2307 731
rect 2309 721 2310 731
rect 2314 721 2315 731
rect 2317 721 2318 731
rect 2350 721 2351 731
rect 2353 721 2354 731
rect 2358 721 2359 731
rect 2361 721 2362 731
rect 2401 721 2402 731
rect 2404 721 2405 731
rect 2541 678 2542 698
rect 2544 678 2545 698
rect 2504 626 2505 646
rect 2507 626 2508 646
rect 2574 631 2575 651
rect 2577 631 2578 651
rect 2617 625 2618 645
rect 2620 625 2621 645
rect 2688 597 2689 637
rect 2691 597 2692 637
rect 2709 597 2710 637
rect 2712 597 2713 637
rect 2734 624 2735 644
rect 2737 624 2738 644
rect 2896 633 2897 693
rect 2899 633 2900 693
rect 2917 633 2918 693
rect 2920 633 2921 693
rect 2938 633 2939 693
rect 2941 633 2942 693
rect 2984 680 2985 700
rect 2987 680 2988 700
rect 3112 666 3113 706
rect 3115 666 3116 706
rect 3133 666 3134 706
rect 3136 666 3137 706
rect 3158 693 3159 713
rect 3161 693 3162 713
rect 3276 658 3277 678
rect 3279 658 3280 678
rect 3297 658 3298 678
rect 3300 658 3301 678
rect 3318 658 3319 678
rect 3321 658 3322 678
rect 3342 660 3343 680
rect 3345 660 3346 680
rect 2270 555 2271 565
rect 2273 555 2274 565
rect 2306 555 2307 565
rect 2309 555 2310 565
rect 2314 555 2315 565
rect 2317 555 2318 565
rect 2350 555 2351 565
rect 2353 555 2354 565
rect 2358 555 2359 565
rect 2361 555 2362 565
rect 2401 555 2402 565
rect 2404 555 2405 565
rect 2270 430 2271 440
rect 2273 430 2274 440
rect 2306 430 2307 440
rect 2309 430 2310 440
rect 2314 430 2315 440
rect 2317 430 2318 440
rect 2350 430 2351 440
rect 2353 430 2354 440
rect 2358 430 2359 440
rect 2361 430 2362 440
rect 2401 430 2402 440
rect 2404 430 2405 440
rect 2556 424 2557 444
rect 2559 424 2560 444
rect 2519 372 2520 392
rect 2522 372 2523 392
rect 2589 377 2590 397
rect 2592 377 2593 397
rect 2632 371 2633 391
rect 2635 371 2636 391
rect 2703 343 2704 383
rect 2706 343 2707 383
rect 2724 343 2725 383
rect 2727 343 2728 383
rect 2749 370 2750 390
rect 2752 370 2753 390
rect 2885 366 2886 446
rect 2888 366 2889 446
rect 2906 366 2907 446
rect 2909 366 2910 446
rect 2927 366 2928 446
rect 2930 366 2931 446
rect 2948 366 2949 446
rect 2951 366 2952 446
rect 2973 433 2974 453
rect 2976 433 2977 453
rect 3072 411 3073 471
rect 3075 411 3076 471
rect 3093 411 3094 471
rect 3096 411 3097 471
rect 3114 411 3115 471
rect 3117 411 3118 471
rect 3160 458 3161 478
rect 3163 458 3164 478
rect 3296 433 3297 473
rect 3299 433 3300 473
rect 3317 433 3318 473
rect 3320 433 3321 473
rect 3342 460 3343 480
rect 3345 460 3346 480
rect 2318 287 2319 297
rect 2321 287 2322 297
rect 2354 287 2355 297
rect 2357 287 2358 297
rect 2362 287 2363 297
rect 2365 287 2366 297
rect 2398 287 2399 297
rect 2401 287 2402 297
rect 2406 287 2407 297
rect 2409 287 2410 297
rect 2449 287 2450 297
rect 2452 287 2453 297
rect 2902 284 2922 285
rect 2902 281 2922 282
rect 2902 263 2922 264
rect 2902 260 2922 261
rect 2902 242 2922 243
rect 2902 239 2922 240
rect 3296 239 3297 259
rect 3299 239 3300 259
rect 2902 221 2922 222
rect 2902 218 2922 219
rect 2909 196 2929 197
rect 2909 193 2929 194
rect 3259 187 3260 207
rect 3262 187 3263 207
rect 3329 192 3330 212
rect 3332 192 3333 212
rect 3372 186 3373 206
rect 3375 186 3376 206
rect 3506 119 3507 129
rect 3509 119 3510 129
rect 3542 119 3543 129
rect 3545 119 3546 129
rect 3550 119 3551 129
rect 3553 119 3554 129
rect 3586 119 3587 129
rect 3589 119 3590 129
rect 3594 119 3595 129
rect 3597 119 3598 129
rect 3637 119 3638 129
rect 3640 119 3641 129
rect 2960 25 2961 35
rect 2963 25 2964 35
rect 2996 25 2997 35
rect 2999 25 3000 35
rect 3004 25 3005 35
rect 3007 25 3008 35
rect 3040 25 3041 35
rect 3043 25 3044 35
rect 3048 25 3049 35
rect 3051 25 3052 35
rect 3091 25 3092 35
rect 3094 25 3095 35
<< pdiffusion >>
rect 2255 1372 2256 1397
rect 2258 1372 2259 1397
rect 2263 1372 2264 1397
rect 2266 1372 2267 1397
rect 2293 1372 2294 1397
rect 2296 1372 2297 1397
rect 2337 1372 2338 1397
rect 2340 1372 2341 1397
rect 2382 1372 2383 1397
rect 2385 1372 2386 1397
rect 2022 1214 2023 1239
rect 2025 1214 2026 1239
rect 2067 1214 2068 1239
rect 2070 1214 2071 1239
rect 2111 1214 2112 1239
rect 2114 1214 2115 1239
rect 2141 1214 2142 1239
rect 2144 1214 2145 1239
rect 2149 1214 2150 1239
rect 2152 1214 2153 1239
rect 2514 1205 2515 1245
rect 2517 1205 2518 1245
rect 2584 1210 2585 1230
rect 2587 1210 2588 1230
rect 2261 1168 2262 1193
rect 2264 1168 2265 1193
rect 2269 1168 2270 1193
rect 2272 1168 2273 1193
rect 2299 1168 2300 1193
rect 2302 1168 2303 1193
rect 2343 1168 2344 1193
rect 2346 1168 2347 1193
rect 2388 1168 2389 1193
rect 2391 1168 2392 1193
rect 2627 1204 2628 1244
rect 2630 1204 2631 1244
rect 2551 1177 2552 1197
rect 2554 1177 2555 1197
rect 2698 1203 2699 1243
rect 2701 1203 2702 1243
rect 2719 1203 2720 1243
rect 2722 1203 2723 1243
rect 2744 1203 2745 1243
rect 2747 1203 2748 1243
rect 2837 1168 2838 1208
rect 2840 1168 2841 1208
rect 2907 1173 2908 1193
rect 2910 1173 2911 1193
rect 2950 1167 2951 1207
rect 2953 1167 2954 1207
rect 3076 1200 3077 1240
rect 3079 1200 3080 1240
rect 3146 1205 3147 1225
rect 3149 1205 3150 1225
rect 3189 1199 3190 1239
rect 3192 1199 3193 1239
rect 2874 1140 2875 1160
rect 2877 1140 2878 1160
rect 3113 1172 3114 1192
rect 3116 1172 3117 1192
rect 3364 1180 3365 1205
rect 3367 1180 3368 1205
rect 3372 1180 3373 1205
rect 3375 1180 3376 1205
rect 3402 1180 3403 1205
rect 3405 1180 3406 1205
rect 3446 1180 3447 1205
rect 3449 1180 3450 1205
rect 3491 1180 3492 1205
rect 3494 1180 3495 1205
rect 2264 1039 2265 1064
rect 2267 1039 2268 1064
rect 2272 1039 2273 1064
rect 2275 1039 2276 1064
rect 2302 1039 2303 1064
rect 2305 1039 2306 1064
rect 2346 1039 2347 1064
rect 2349 1039 2350 1064
rect 2391 1039 2392 1064
rect 2394 1039 2395 1064
rect 3367 1044 3368 1069
rect 3370 1044 3371 1069
rect 3375 1044 3376 1069
rect 3378 1044 3379 1069
rect 3405 1044 3406 1069
rect 3408 1044 3409 1069
rect 3449 1044 3450 1069
rect 3452 1044 3453 1069
rect 3494 1044 3495 1069
rect 3497 1044 3498 1069
rect 2494 911 2495 951
rect 2497 911 2498 951
rect 2564 916 2565 936
rect 2567 916 2568 936
rect 2274 878 2275 903
rect 2277 878 2278 903
rect 2282 878 2283 903
rect 2285 878 2286 903
rect 2312 878 2313 903
rect 2315 878 2316 903
rect 2356 878 2357 903
rect 2359 878 2360 903
rect 2401 878 2402 903
rect 2404 878 2405 903
rect 2607 910 2608 950
rect 2610 910 2611 950
rect 2531 883 2532 903
rect 2534 883 2535 903
rect 2678 909 2679 949
rect 2681 909 2682 949
rect 2699 909 2700 949
rect 2702 909 2703 949
rect 2724 909 2725 949
rect 2727 909 2728 949
rect 2914 943 2915 983
rect 2917 943 2918 983
rect 2935 943 2936 983
rect 2938 943 2939 983
rect 2960 943 2961 983
rect 2963 943 2964 983
rect 3030 910 3031 990
rect 3033 910 3034 990
rect 3051 910 3052 990
rect 3054 910 3055 990
rect 3076 910 3077 950
rect 3079 910 3080 950
rect 2274 753 2275 778
rect 2277 753 2278 778
rect 2282 753 2283 778
rect 2285 753 2286 778
rect 2312 753 2313 778
rect 2315 753 2316 778
rect 2356 753 2357 778
rect 2359 753 2360 778
rect 2401 753 2402 778
rect 2404 753 2405 778
rect 2504 666 2505 706
rect 2507 666 2508 706
rect 2574 671 2575 691
rect 2577 671 2578 691
rect 2617 665 2618 705
rect 2620 665 2621 705
rect 2896 720 2897 760
rect 2899 720 2900 760
rect 2917 720 2918 760
rect 2920 720 2921 760
rect 2938 720 2939 760
rect 2941 720 2942 760
rect 2984 720 2985 760
rect 2987 720 2988 760
rect 3112 733 3113 773
rect 3115 733 3116 773
rect 3133 733 3134 773
rect 3136 733 3137 773
rect 3158 733 3159 773
rect 3161 733 3162 773
rect 2541 638 2542 658
rect 2544 638 2545 658
rect 2688 664 2689 704
rect 2691 664 2692 704
rect 2709 664 2710 704
rect 2712 664 2713 704
rect 2734 664 2735 704
rect 2737 664 2738 704
rect 2274 587 2275 612
rect 2277 587 2278 612
rect 2282 587 2283 612
rect 2285 587 2286 612
rect 2312 587 2313 612
rect 2315 587 2316 612
rect 2356 587 2357 612
rect 2359 587 2360 612
rect 2401 587 2402 612
rect 2404 587 2405 612
rect 3276 699 3277 819
rect 3279 699 3280 819
rect 3297 699 3298 819
rect 3300 699 3301 819
rect 3318 699 3319 819
rect 3321 699 3322 819
rect 3342 700 3343 740
rect 3345 700 3346 740
rect 2274 462 2275 487
rect 2277 462 2278 487
rect 2282 462 2283 487
rect 2285 462 2286 487
rect 2312 462 2313 487
rect 2315 462 2316 487
rect 2356 462 2357 487
rect 2359 462 2360 487
rect 2401 462 2402 487
rect 2404 462 2405 487
rect 2885 473 2886 513
rect 2888 473 2889 513
rect 2906 473 2907 513
rect 2909 473 2910 513
rect 2927 473 2928 513
rect 2930 473 2931 513
rect 2948 473 2949 513
rect 2951 473 2952 513
rect 2973 473 2974 513
rect 2976 473 2977 513
rect 3072 498 3073 538
rect 3075 498 3076 538
rect 3093 498 3094 538
rect 3096 498 3097 538
rect 3114 498 3115 538
rect 3117 498 3118 538
rect 3160 498 3161 538
rect 3163 498 3164 538
rect 3296 500 3297 540
rect 3299 500 3300 540
rect 3317 500 3318 540
rect 3320 500 3321 540
rect 3342 500 3343 540
rect 3345 500 3346 540
rect 2519 412 2520 452
rect 2522 412 2523 452
rect 2589 417 2590 437
rect 2592 417 2593 437
rect 2632 411 2633 451
rect 2635 411 2636 451
rect 2556 384 2557 404
rect 2559 384 2560 404
rect 2703 410 2704 450
rect 2706 410 2707 450
rect 2724 410 2725 450
rect 2727 410 2728 450
rect 2749 410 2750 450
rect 2752 410 2753 450
rect 2322 319 2323 344
rect 2325 319 2326 344
rect 2330 319 2331 344
rect 2333 319 2334 344
rect 2360 319 2361 344
rect 2363 319 2364 344
rect 2404 319 2405 344
rect 2407 319 2408 344
rect 2449 319 2450 344
rect 2452 319 2453 344
rect 2949 284 3109 285
rect 2949 281 3109 282
rect 2949 263 3109 264
rect 2949 260 3109 261
rect 2949 242 3109 243
rect 2949 239 3109 240
rect 3259 227 3260 267
rect 3262 227 3263 267
rect 3329 232 3330 252
rect 3332 232 3333 252
rect 2949 221 3109 222
rect 2949 218 3109 219
rect 3372 226 3373 266
rect 3375 226 3376 266
rect 2949 196 2989 197
rect 2949 193 2989 194
rect 3296 199 3297 219
rect 3299 199 3300 219
rect 3510 151 3511 176
rect 3513 151 3514 176
rect 3518 151 3519 176
rect 3521 151 3522 176
rect 3548 151 3549 176
rect 3551 151 3552 176
rect 3592 151 3593 176
rect 3595 151 3596 176
rect 3637 151 3638 176
rect 3640 151 3641 176
rect 2964 57 2965 82
rect 2967 57 2968 82
rect 2972 57 2973 82
rect 2975 57 2976 82
rect 3002 57 3003 82
rect 3005 57 3006 82
rect 3046 57 3047 82
rect 3049 57 3050 82
rect 3091 57 3092 82
rect 3094 57 3095 82
<< ndcontact >>
rect 2247 1340 2251 1350
rect 2255 1340 2259 1350
rect 2283 1340 2287 1350
rect 2291 1340 2295 1350
rect 2299 1340 2303 1350
rect 2327 1340 2331 1350
rect 2335 1340 2339 1350
rect 2343 1340 2347 1350
rect 2378 1340 2382 1350
rect 2386 1340 2390 1350
rect 2018 1261 2022 1271
rect 2026 1261 2030 1271
rect 2061 1261 2065 1271
rect 2069 1261 2073 1271
rect 2077 1261 2081 1271
rect 2105 1261 2109 1271
rect 2113 1261 2117 1271
rect 2121 1261 2125 1271
rect 2149 1261 2153 1271
rect 2157 1261 2161 1271
rect 2547 1217 2551 1237
rect 2555 1217 2559 1237
rect 2510 1165 2514 1185
rect 2518 1165 2522 1185
rect 2580 1170 2584 1190
rect 2588 1170 2592 1190
rect 2623 1164 2627 1184
rect 2631 1164 2635 1184
rect 2253 1136 2257 1146
rect 2261 1136 2265 1146
rect 2289 1136 2293 1146
rect 2297 1136 2301 1146
rect 2305 1136 2309 1146
rect 2333 1136 2337 1146
rect 2341 1136 2345 1146
rect 2349 1136 2353 1146
rect 2384 1136 2388 1146
rect 2392 1136 2396 1146
rect 2694 1136 2698 1176
rect 2702 1136 2719 1176
rect 2723 1136 2727 1176
rect 2740 1163 2744 1183
rect 2748 1163 2752 1183
rect 2870 1180 2874 1200
rect 2878 1180 2882 1200
rect 3109 1212 3113 1232
rect 3117 1212 3121 1232
rect 2833 1128 2837 1148
rect 2841 1128 2845 1148
rect 2903 1133 2907 1153
rect 2911 1133 2915 1153
rect 3072 1160 3076 1180
rect 3080 1160 3084 1180
rect 3142 1165 3146 1185
rect 3150 1165 3154 1185
rect 3185 1159 3189 1179
rect 3193 1159 3197 1179
rect 3356 1148 3360 1158
rect 3364 1148 3368 1158
rect 3392 1148 3396 1158
rect 3400 1148 3404 1158
rect 3408 1148 3412 1158
rect 3436 1148 3440 1158
rect 3444 1148 3448 1158
rect 3452 1148 3456 1158
rect 3487 1148 3491 1158
rect 3495 1148 3499 1158
rect 2946 1127 2950 1147
rect 2954 1127 2958 1147
rect 2256 1007 2260 1017
rect 2264 1007 2268 1017
rect 2292 1007 2296 1017
rect 2300 1007 2304 1017
rect 2308 1007 2312 1017
rect 2336 1007 2340 1017
rect 2344 1007 2348 1017
rect 2352 1007 2356 1017
rect 2387 1007 2391 1017
rect 2395 1007 2399 1017
rect 3359 1012 3363 1022
rect 3367 1012 3371 1022
rect 3395 1012 3399 1022
rect 3403 1012 3407 1022
rect 3411 1012 3415 1022
rect 3439 1012 3443 1022
rect 3447 1012 3451 1022
rect 3455 1012 3459 1022
rect 3490 1012 3494 1022
rect 3498 1012 3502 1022
rect 2527 923 2531 943
rect 2535 923 2539 943
rect 2490 871 2494 891
rect 2498 871 2502 891
rect 2560 876 2564 896
rect 2568 876 2572 896
rect 2603 870 2607 890
rect 2611 870 2615 890
rect 2266 846 2270 856
rect 2274 846 2278 856
rect 2302 846 2306 856
rect 2310 846 2314 856
rect 2318 846 2322 856
rect 2346 846 2350 856
rect 2354 846 2358 856
rect 2362 846 2366 856
rect 2397 846 2401 856
rect 2405 846 2409 856
rect 2674 842 2678 882
rect 2682 842 2699 882
rect 2703 842 2707 882
rect 2720 869 2724 889
rect 2728 869 2732 889
rect 2910 876 2914 916
rect 2918 876 2935 916
rect 2939 876 2943 916
rect 2956 903 2960 923
rect 2964 903 2968 923
rect 3026 868 3030 888
rect 3034 868 3038 888
rect 3047 868 3051 888
rect 3055 868 3059 888
rect 3072 870 3076 890
rect 3080 870 3084 890
rect 2266 721 2270 731
rect 2274 721 2278 731
rect 2302 721 2306 731
rect 2310 721 2314 731
rect 2318 721 2322 731
rect 2346 721 2350 731
rect 2354 721 2358 731
rect 2362 721 2366 731
rect 2397 721 2401 731
rect 2405 721 2409 731
rect 2537 678 2541 698
rect 2545 678 2549 698
rect 2500 626 2504 646
rect 2508 626 2512 646
rect 2570 631 2574 651
rect 2578 631 2582 651
rect 2613 625 2617 645
rect 2621 625 2625 645
rect 2684 597 2688 637
rect 2692 597 2709 637
rect 2713 597 2717 637
rect 2730 624 2734 644
rect 2738 624 2742 644
rect 2892 633 2896 693
rect 2900 633 2904 693
rect 2913 633 2917 693
rect 2921 633 2925 693
rect 2934 633 2938 693
rect 2942 633 2946 693
rect 2980 680 2984 700
rect 2988 680 2992 700
rect 3108 666 3112 706
rect 3116 666 3133 706
rect 3137 666 3141 706
rect 3154 693 3158 713
rect 3162 693 3166 713
rect 3272 658 3276 678
rect 3280 658 3284 678
rect 3293 658 3297 678
rect 3301 658 3305 678
rect 3314 658 3318 678
rect 3322 658 3326 678
rect 3338 660 3342 680
rect 3346 660 3350 680
rect 2266 555 2270 565
rect 2274 555 2278 565
rect 2302 555 2306 565
rect 2310 555 2314 565
rect 2318 555 2322 565
rect 2346 555 2350 565
rect 2354 555 2358 565
rect 2362 555 2366 565
rect 2397 555 2401 565
rect 2405 555 2409 565
rect 2266 430 2270 440
rect 2274 430 2278 440
rect 2302 430 2306 440
rect 2310 430 2314 440
rect 2318 430 2322 440
rect 2346 430 2350 440
rect 2354 430 2358 440
rect 2362 430 2366 440
rect 2397 430 2401 440
rect 2405 430 2409 440
rect 2552 424 2556 444
rect 2560 424 2564 444
rect 2515 372 2519 392
rect 2523 372 2527 392
rect 2585 377 2589 397
rect 2593 377 2597 397
rect 2628 371 2632 391
rect 2636 371 2640 391
rect 2699 343 2703 383
rect 2707 343 2724 383
rect 2728 343 2732 383
rect 2745 370 2749 390
rect 2753 370 2757 390
rect 2881 366 2885 446
rect 2889 366 2893 446
rect 2902 366 2906 446
rect 2910 366 2914 446
rect 2923 366 2927 446
rect 2931 366 2935 446
rect 2944 366 2948 446
rect 2952 366 2956 446
rect 2969 433 2973 453
rect 2977 433 2981 453
rect 3068 411 3072 471
rect 3076 411 3080 471
rect 3089 411 3093 471
rect 3097 411 3101 471
rect 3110 411 3114 471
rect 3118 411 3122 471
rect 3156 458 3160 478
rect 3164 458 3168 478
rect 3292 433 3296 473
rect 3300 433 3317 473
rect 3321 433 3325 473
rect 3338 460 3342 480
rect 3346 460 3350 480
rect 2314 287 2318 297
rect 2322 287 2326 297
rect 2350 287 2354 297
rect 2358 287 2362 297
rect 2366 287 2370 297
rect 2394 287 2398 297
rect 2402 287 2406 297
rect 2410 287 2414 297
rect 2445 287 2449 297
rect 2453 287 2457 297
rect 2902 285 2922 289
rect 2902 277 2922 281
rect 2902 264 2922 268
rect 2902 256 2922 260
rect 2902 243 2922 247
rect 2902 235 2922 239
rect 3292 239 3296 259
rect 3300 239 3304 259
rect 2902 222 2922 226
rect 2902 214 2922 218
rect 2909 197 2929 201
rect 2909 189 2929 193
rect 3255 187 3259 207
rect 3263 187 3267 207
rect 3325 192 3329 212
rect 3333 192 3337 212
rect 3368 186 3372 206
rect 3376 186 3380 206
rect 3502 119 3506 129
rect 3510 119 3514 129
rect 3538 119 3542 129
rect 3546 119 3550 129
rect 3554 119 3558 129
rect 3582 119 3586 129
rect 3590 119 3594 129
rect 3598 119 3602 129
rect 3633 119 3637 129
rect 3641 119 3645 129
rect 2956 25 2960 35
rect 2964 25 2968 35
rect 2992 25 2996 35
rect 3000 25 3004 35
rect 3008 25 3012 35
rect 3036 25 3040 35
rect 3044 25 3048 35
rect 3052 25 3056 35
rect 3087 25 3091 35
rect 3095 25 3099 35
<< pdcontact >>
rect 2251 1372 2255 1397
rect 2259 1372 2263 1397
rect 2267 1372 2271 1397
rect 2289 1372 2293 1397
rect 2297 1372 2301 1397
rect 2333 1372 2337 1397
rect 2341 1372 2345 1397
rect 2378 1372 2382 1397
rect 2386 1372 2390 1397
rect 2018 1214 2022 1239
rect 2026 1214 2030 1239
rect 2063 1214 2067 1239
rect 2071 1214 2075 1239
rect 2107 1214 2111 1239
rect 2115 1214 2119 1239
rect 2137 1214 2141 1239
rect 2145 1214 2149 1239
rect 2153 1214 2157 1239
rect 2510 1205 2514 1245
rect 2518 1205 2522 1245
rect 2580 1210 2584 1230
rect 2588 1210 2592 1230
rect 2257 1168 2261 1193
rect 2265 1168 2269 1193
rect 2273 1168 2277 1193
rect 2295 1168 2299 1193
rect 2303 1168 2307 1193
rect 2339 1168 2343 1193
rect 2347 1168 2351 1193
rect 2384 1168 2388 1193
rect 2392 1168 2396 1193
rect 2623 1204 2627 1244
rect 2631 1204 2635 1244
rect 2547 1177 2551 1197
rect 2555 1177 2559 1197
rect 2694 1203 2698 1243
rect 2702 1203 2719 1243
rect 2723 1203 2727 1243
rect 2740 1203 2744 1243
rect 2748 1203 2752 1243
rect 2833 1168 2837 1208
rect 2841 1168 2845 1208
rect 2903 1173 2907 1193
rect 2911 1173 2915 1193
rect 2946 1167 2950 1207
rect 2954 1167 2958 1207
rect 3072 1200 3076 1240
rect 3080 1200 3084 1240
rect 3142 1205 3146 1225
rect 3150 1205 3154 1225
rect 3185 1199 3189 1239
rect 3193 1199 3197 1239
rect 2870 1140 2874 1160
rect 2878 1140 2882 1160
rect 3109 1172 3113 1192
rect 3117 1172 3121 1192
rect 3360 1180 3364 1205
rect 3368 1180 3372 1205
rect 3376 1180 3380 1205
rect 3398 1180 3402 1205
rect 3406 1180 3410 1205
rect 3442 1180 3446 1205
rect 3450 1180 3454 1205
rect 3487 1180 3491 1205
rect 3495 1180 3499 1205
rect 2260 1039 2264 1064
rect 2268 1039 2272 1064
rect 2276 1039 2280 1064
rect 2298 1039 2302 1064
rect 2306 1039 2310 1064
rect 2342 1039 2346 1064
rect 2350 1039 2354 1064
rect 2387 1039 2391 1064
rect 2395 1039 2399 1064
rect 3363 1044 3367 1069
rect 3371 1044 3375 1069
rect 3379 1044 3383 1069
rect 3401 1044 3405 1069
rect 3409 1044 3413 1069
rect 3445 1044 3449 1069
rect 3453 1044 3457 1069
rect 3490 1044 3494 1069
rect 3498 1044 3502 1069
rect 2490 911 2494 951
rect 2498 911 2502 951
rect 2560 916 2564 936
rect 2568 916 2572 936
rect 2270 878 2274 903
rect 2278 878 2282 903
rect 2286 878 2290 903
rect 2308 878 2312 903
rect 2316 878 2320 903
rect 2352 878 2356 903
rect 2360 878 2364 903
rect 2397 878 2401 903
rect 2405 878 2409 903
rect 2603 910 2607 950
rect 2611 910 2615 950
rect 2527 883 2531 903
rect 2535 883 2539 903
rect 2674 909 2678 949
rect 2682 909 2699 949
rect 2703 909 2707 949
rect 2720 909 2724 949
rect 2728 909 2732 949
rect 2910 943 2914 983
rect 2918 943 2935 983
rect 2939 943 2943 983
rect 2956 943 2960 983
rect 2964 943 2968 983
rect 3026 910 3030 990
rect 3034 910 3038 990
rect 3047 910 3051 990
rect 3055 910 3059 990
rect 3072 910 3076 950
rect 3080 910 3084 950
rect 2270 753 2274 778
rect 2278 753 2282 778
rect 2286 753 2290 778
rect 2308 753 2312 778
rect 2316 753 2320 778
rect 2352 753 2356 778
rect 2360 753 2364 778
rect 2397 753 2401 778
rect 2405 753 2409 778
rect 2500 666 2504 706
rect 2508 666 2512 706
rect 2570 671 2574 691
rect 2578 671 2582 691
rect 2613 665 2617 705
rect 2621 665 2625 705
rect 2892 720 2896 760
rect 2900 720 2917 760
rect 2921 720 2938 760
rect 2942 720 2946 760
rect 2980 720 2984 760
rect 2988 720 2992 760
rect 3108 733 3112 773
rect 3116 733 3133 773
rect 3137 733 3141 773
rect 3154 733 3158 773
rect 3162 733 3166 773
rect 2537 638 2541 658
rect 2545 638 2549 658
rect 2684 664 2688 704
rect 2692 664 2709 704
rect 2713 664 2717 704
rect 2730 664 2734 704
rect 2738 664 2742 704
rect 2270 587 2274 612
rect 2278 587 2282 612
rect 2286 587 2290 612
rect 2308 587 2312 612
rect 2316 587 2320 612
rect 2352 587 2356 612
rect 2360 587 2364 612
rect 2397 587 2401 612
rect 2405 587 2409 612
rect 3272 699 3276 819
rect 3280 699 3284 819
rect 3293 699 3297 819
rect 3301 699 3305 819
rect 3314 699 3318 819
rect 3322 699 3326 819
rect 3338 700 3342 740
rect 3346 700 3350 740
rect 2270 462 2274 487
rect 2278 462 2282 487
rect 2286 462 2290 487
rect 2308 462 2312 487
rect 2316 462 2320 487
rect 2352 462 2356 487
rect 2360 462 2364 487
rect 2397 462 2401 487
rect 2405 462 2409 487
rect 2881 473 2885 513
rect 2889 473 2906 513
rect 2910 473 2927 513
rect 2931 473 2948 513
rect 2952 473 2956 513
rect 2969 473 2973 513
rect 2977 473 2981 513
rect 3068 498 3072 538
rect 3076 498 3093 538
rect 3097 498 3114 538
rect 3118 498 3122 538
rect 3156 498 3160 538
rect 3164 498 3168 538
rect 3292 500 3296 540
rect 3300 500 3317 540
rect 3321 500 3325 540
rect 3338 500 3342 540
rect 3346 500 3350 540
rect 2515 412 2519 452
rect 2523 412 2527 452
rect 2585 417 2589 437
rect 2593 417 2597 437
rect 2628 411 2632 451
rect 2636 411 2640 451
rect 2552 384 2556 404
rect 2560 384 2564 404
rect 2699 410 2703 450
rect 2707 410 2724 450
rect 2728 410 2732 450
rect 2745 410 2749 450
rect 2753 410 2757 450
rect 2318 319 2322 344
rect 2326 319 2330 344
rect 2334 319 2338 344
rect 2356 319 2360 344
rect 2364 319 2368 344
rect 2400 319 2404 344
rect 2408 319 2412 344
rect 2445 319 2449 344
rect 2453 319 2457 344
rect 2949 285 3109 289
rect 2949 277 3109 281
rect 2949 264 3109 268
rect 2949 256 3109 260
rect 2949 243 3109 247
rect 2949 235 3109 239
rect 3255 227 3259 267
rect 3263 227 3267 267
rect 3325 232 3329 252
rect 3333 232 3337 252
rect 2949 222 3109 226
rect 2949 214 3109 218
rect 3368 226 3372 266
rect 3376 226 3380 266
rect 2949 197 2989 201
rect 2949 189 2989 193
rect 3292 199 3296 219
rect 3300 199 3304 219
rect 3506 151 3510 176
rect 3514 151 3518 176
rect 3522 151 3526 176
rect 3544 151 3548 176
rect 3552 151 3556 176
rect 3588 151 3592 176
rect 3596 151 3600 176
rect 3633 151 3637 176
rect 3641 151 3645 176
rect 2960 57 2964 82
rect 2968 57 2972 82
rect 2976 57 2980 82
rect 2998 57 3002 82
rect 3006 57 3010 82
rect 3042 57 3046 82
rect 3050 57 3054 82
rect 3087 57 3091 82
rect 3095 57 3099 82
<< polysilicon >>
rect 2256 1397 2258 1400
rect 2264 1397 2266 1400
rect 2294 1397 2296 1400
rect 2338 1397 2340 1400
rect 2383 1397 2385 1400
rect 2256 1365 2258 1372
rect 2251 1361 2258 1365
rect 2252 1350 2254 1361
rect 2264 1353 2266 1372
rect 2294 1364 2296 1372
rect 2338 1364 2340 1372
rect 2288 1362 2296 1364
rect 2332 1362 2340 1364
rect 2288 1350 2290 1362
rect 2296 1350 2298 1359
rect 2332 1350 2334 1362
rect 2340 1350 2342 1359
rect 2383 1350 2385 1372
rect 2252 1337 2254 1340
rect 2288 1337 2290 1340
rect 2296 1337 2298 1340
rect 2332 1337 2334 1340
rect 2340 1337 2342 1340
rect 2383 1337 2385 1340
rect 2023 1271 2025 1274
rect 2066 1271 2068 1274
rect 2074 1271 2076 1274
rect 2110 1271 2112 1274
rect 2118 1271 2120 1274
rect 2154 1271 2156 1274
rect 2023 1239 2025 1261
rect 2066 1252 2068 1261
rect 2074 1249 2076 1261
rect 2110 1252 2112 1261
rect 2118 1249 2120 1261
rect 2068 1247 2076 1249
rect 2112 1247 2120 1249
rect 2068 1239 2070 1247
rect 2112 1239 2114 1247
rect 2142 1239 2144 1258
rect 2154 1250 2156 1261
rect 2150 1246 2157 1250
rect 2150 1239 2152 1246
rect 2515 1245 2517 1249
rect 2023 1211 2025 1214
rect 2068 1211 2070 1214
rect 2112 1211 2114 1214
rect 2142 1211 2144 1214
rect 2150 1211 2152 1214
rect 2628 1244 2630 1248
rect 2552 1237 2554 1244
rect 2585 1230 2587 1244
rect 2552 1214 2554 1217
rect 2585 1207 2587 1210
rect 2262 1193 2264 1196
rect 2270 1193 2272 1196
rect 2300 1193 2302 1196
rect 2344 1193 2346 1196
rect 2389 1193 2391 1196
rect 2515 1185 2517 1205
rect 2699 1243 2701 1247
rect 2720 1243 2722 1262
rect 2745 1243 2747 1247
rect 2552 1197 2554 1200
rect 2262 1161 2264 1168
rect 2257 1157 2264 1161
rect 2258 1146 2260 1157
rect 2270 1149 2272 1168
rect 2300 1160 2302 1168
rect 2344 1160 2346 1168
rect 2294 1158 2302 1160
rect 2338 1158 2346 1160
rect 2294 1146 2296 1158
rect 2302 1146 2304 1155
rect 2338 1146 2340 1158
rect 2346 1146 2348 1155
rect 2389 1146 2391 1168
rect 2585 1190 2587 1193
rect 2515 1162 2517 1165
rect 2552 1163 2554 1177
rect 2628 1184 2630 1204
rect 3077 1240 3079 1244
rect 2838 1208 2840 1212
rect 2585 1163 2587 1170
rect 2699 1176 2701 1203
rect 2720 1176 2722 1203
rect 2745 1183 2747 1203
rect 2628 1161 2630 1164
rect 2951 1207 2953 1211
rect 2875 1200 2877 1207
rect 2908 1193 2910 1207
rect 2875 1177 2877 1180
rect 2908 1170 2910 1173
rect 2745 1160 2747 1163
rect 2838 1148 2840 1168
rect 3190 1239 3192 1243
rect 3114 1232 3116 1239
rect 3147 1225 3149 1239
rect 3114 1209 3116 1212
rect 3147 1202 3149 1205
rect 3077 1180 3079 1200
rect 3365 1205 3367 1208
rect 3373 1205 3375 1208
rect 3403 1205 3405 1208
rect 3447 1205 3449 1208
rect 3492 1205 3494 1208
rect 3114 1192 3116 1195
rect 2875 1160 2877 1163
rect 2258 1133 2260 1136
rect 2294 1133 2296 1136
rect 2302 1133 2304 1136
rect 2338 1133 2340 1136
rect 2346 1133 2348 1136
rect 2389 1133 2391 1136
rect 2699 1133 2701 1136
rect 2720 1133 2722 1136
rect 2908 1153 2910 1156
rect 2838 1125 2840 1128
rect 2875 1126 2877 1140
rect 2951 1147 2953 1167
rect 3147 1185 3149 1188
rect 3077 1157 3079 1160
rect 3114 1158 3116 1172
rect 3190 1179 3192 1199
rect 3147 1158 3149 1165
rect 3365 1173 3367 1180
rect 3360 1169 3367 1173
rect 3190 1156 3192 1159
rect 3361 1158 3363 1169
rect 3373 1161 3375 1180
rect 3403 1172 3405 1180
rect 3447 1172 3449 1180
rect 3397 1170 3405 1172
rect 3441 1170 3449 1172
rect 3397 1158 3399 1170
rect 3405 1158 3407 1167
rect 3441 1158 3443 1170
rect 3449 1158 3451 1167
rect 3492 1158 3494 1180
rect 2908 1126 2910 1133
rect 3361 1145 3363 1148
rect 3397 1145 3399 1148
rect 3405 1145 3407 1148
rect 3441 1145 3443 1148
rect 3449 1145 3451 1148
rect 3492 1145 3494 1148
rect 2951 1124 2953 1127
rect 3368 1069 3370 1072
rect 3376 1069 3378 1072
rect 3406 1069 3408 1072
rect 3450 1069 3452 1072
rect 3495 1069 3497 1072
rect 2265 1064 2267 1067
rect 2273 1064 2275 1067
rect 2303 1064 2305 1067
rect 2347 1064 2349 1067
rect 2392 1064 2394 1067
rect 2265 1032 2267 1039
rect 2260 1028 2267 1032
rect 2261 1017 2263 1028
rect 2273 1020 2275 1039
rect 2303 1031 2305 1039
rect 2347 1031 2349 1039
rect 2297 1029 2305 1031
rect 2341 1029 2349 1031
rect 2297 1017 2299 1029
rect 2305 1017 2307 1026
rect 2341 1017 2343 1029
rect 2349 1017 2351 1026
rect 2392 1017 2394 1039
rect 3368 1037 3370 1044
rect 3363 1033 3370 1037
rect 3364 1022 3366 1033
rect 3376 1025 3378 1044
rect 3406 1036 3408 1044
rect 3450 1036 3452 1044
rect 3400 1034 3408 1036
rect 3444 1034 3452 1036
rect 3400 1022 3402 1034
rect 3408 1022 3410 1031
rect 3444 1022 3446 1034
rect 3452 1022 3454 1031
rect 3495 1022 3497 1044
rect 3364 1009 3366 1012
rect 3400 1009 3402 1012
rect 3408 1009 3410 1012
rect 3444 1009 3446 1012
rect 3452 1009 3454 1012
rect 3495 1009 3497 1012
rect 2261 1004 2263 1007
rect 2297 1004 2299 1007
rect 2305 1004 2307 1007
rect 2341 1004 2343 1007
rect 2349 1004 2351 1007
rect 2392 1004 2394 1007
rect 2915 983 2917 987
rect 2936 983 2938 1002
rect 3031 990 3033 993
rect 3052 990 3054 1007
rect 2961 983 2963 987
rect 2495 951 2497 955
rect 2608 950 2610 954
rect 2532 943 2534 950
rect 2565 936 2567 950
rect 2532 920 2534 923
rect 2565 913 2567 916
rect 2275 903 2277 906
rect 2283 903 2285 906
rect 2313 903 2315 906
rect 2357 903 2359 906
rect 2402 903 2404 906
rect 2495 891 2497 911
rect 2679 949 2681 953
rect 2700 949 2702 968
rect 2725 949 2727 953
rect 2532 903 2534 906
rect 2275 871 2277 878
rect 2270 867 2277 871
rect 2271 856 2273 867
rect 2283 859 2285 878
rect 2313 870 2315 878
rect 2357 870 2359 878
rect 2307 868 2315 870
rect 2351 868 2359 870
rect 2307 856 2309 868
rect 2315 856 2317 865
rect 2351 856 2353 868
rect 2359 856 2361 865
rect 2402 856 2404 878
rect 2565 896 2567 899
rect 2495 868 2497 871
rect 2532 869 2534 883
rect 2608 890 2610 910
rect 2915 916 2917 943
rect 2936 916 2938 943
rect 2961 923 2963 943
rect 2565 869 2567 876
rect 2679 882 2681 909
rect 2700 882 2702 909
rect 2725 889 2727 909
rect 2608 867 2610 870
rect 2271 843 2273 846
rect 2307 843 2309 846
rect 2315 843 2317 846
rect 2351 843 2353 846
rect 2359 843 2361 846
rect 2402 843 2404 846
rect 3077 950 3079 954
rect 2961 900 2963 903
rect 3031 888 3033 910
rect 3052 888 3054 910
rect 3077 890 3079 910
rect 2915 873 2917 876
rect 2936 873 2938 876
rect 2725 866 2727 869
rect 3031 865 3033 868
rect 3052 865 3054 868
rect 3077 867 3079 870
rect 2679 839 2681 842
rect 2700 839 2702 842
rect 3277 819 3279 827
rect 3298 819 3300 841
rect 3319 819 3321 851
rect 2275 778 2277 781
rect 2283 778 2285 781
rect 2313 778 2315 781
rect 2357 778 2359 781
rect 2402 778 2404 781
rect 2897 760 2899 764
rect 2918 760 2920 779
rect 2939 760 2941 792
rect 3113 773 3115 777
rect 3134 773 3136 792
rect 3159 773 3161 777
rect 2985 760 2987 764
rect 2275 746 2277 753
rect 2270 742 2277 746
rect 2271 731 2273 742
rect 2283 734 2285 753
rect 2313 745 2315 753
rect 2357 745 2359 753
rect 2307 743 2315 745
rect 2351 743 2359 745
rect 2307 731 2309 743
rect 2315 731 2317 740
rect 2351 731 2353 743
rect 2359 731 2361 740
rect 2402 731 2404 753
rect 2271 718 2273 721
rect 2307 718 2309 721
rect 2315 718 2317 721
rect 2351 718 2353 721
rect 2359 718 2361 721
rect 2402 718 2404 721
rect 2505 706 2507 710
rect 2618 705 2620 709
rect 2542 698 2544 705
rect 2575 691 2577 705
rect 2542 675 2544 678
rect 2575 668 2577 671
rect 2505 646 2507 666
rect 2689 704 2691 708
rect 2710 704 2712 723
rect 2735 704 2737 708
rect 2542 658 2544 661
rect 2575 651 2577 654
rect 2505 623 2507 626
rect 2542 624 2544 638
rect 2618 645 2620 665
rect 2897 693 2899 720
rect 2918 693 2920 720
rect 2939 693 2941 720
rect 2985 700 2987 720
rect 3113 706 3115 733
rect 3134 706 3136 733
rect 3159 713 3161 733
rect 2575 624 2577 631
rect 2689 637 2691 664
rect 2710 637 2712 664
rect 2735 644 2737 664
rect 2618 622 2620 625
rect 2275 612 2277 615
rect 2283 612 2285 615
rect 2313 612 2315 615
rect 2357 612 2359 615
rect 2402 612 2404 615
rect 2985 677 2987 680
rect 3343 740 3345 744
rect 3159 690 3161 693
rect 3277 678 3279 699
rect 3298 678 3300 699
rect 3319 678 3321 699
rect 3343 680 3345 700
rect 3113 663 3115 666
rect 3134 663 3136 666
rect 3277 655 3279 658
rect 3298 655 3300 658
rect 3319 655 3321 658
rect 3343 657 3345 660
rect 2897 629 2899 633
rect 2918 629 2920 633
rect 2939 629 2941 633
rect 2735 621 2737 624
rect 2689 594 2691 597
rect 2710 594 2712 597
rect 2275 580 2277 587
rect 2270 576 2277 580
rect 2271 565 2273 576
rect 2283 568 2285 587
rect 2313 579 2315 587
rect 2357 579 2359 587
rect 2307 577 2315 579
rect 2351 577 2359 579
rect 2307 565 2309 577
rect 2315 565 2317 574
rect 2351 565 2353 577
rect 2359 565 2361 574
rect 2402 565 2404 587
rect 2271 552 2273 555
rect 2307 552 2309 555
rect 2315 552 2317 555
rect 2351 552 2353 555
rect 2359 552 2361 555
rect 2402 552 2404 555
rect 2886 513 2888 517
rect 2907 513 2909 532
rect 2928 513 2930 559
rect 2949 513 2951 570
rect 3073 538 3075 542
rect 3094 538 3096 559
rect 3115 538 3117 570
rect 3161 538 3163 542
rect 3297 540 3299 544
rect 3318 540 3320 559
rect 3343 540 3345 544
rect 2974 513 2976 517
rect 2275 487 2277 490
rect 2283 487 2285 490
rect 2313 487 2315 490
rect 2357 487 2359 490
rect 2402 487 2404 490
rect 2275 455 2277 462
rect 2270 451 2277 455
rect 2271 440 2273 451
rect 2283 443 2285 462
rect 2313 454 2315 462
rect 2357 454 2359 462
rect 2307 452 2315 454
rect 2351 452 2359 454
rect 2307 440 2309 452
rect 2315 440 2317 449
rect 2351 440 2353 452
rect 2359 440 2361 449
rect 2402 440 2404 462
rect 2520 452 2522 456
rect 2271 427 2273 430
rect 2307 427 2309 430
rect 2315 427 2317 430
rect 2351 427 2353 430
rect 2359 427 2361 430
rect 2402 427 2404 430
rect 2633 451 2635 455
rect 2557 444 2559 451
rect 2590 437 2592 451
rect 2557 421 2559 424
rect 2590 414 2592 417
rect 2520 392 2522 412
rect 2704 450 2706 454
rect 2725 450 2727 469
rect 2750 450 2752 454
rect 2557 404 2559 407
rect 2590 397 2592 400
rect 2520 369 2522 372
rect 2557 370 2559 384
rect 2633 391 2635 411
rect 2886 446 2888 473
rect 2907 446 2909 473
rect 2928 446 2930 473
rect 2949 446 2951 473
rect 2974 453 2976 473
rect 3073 471 3075 498
rect 3094 471 3096 498
rect 3115 471 3117 498
rect 3161 478 3163 498
rect 2590 370 2592 377
rect 2704 383 2706 410
rect 2725 383 2727 410
rect 2750 390 2752 410
rect 2633 368 2635 371
rect 2323 344 2325 347
rect 2331 344 2333 347
rect 2361 344 2363 347
rect 2405 344 2407 347
rect 2450 344 2452 347
rect 2750 367 2752 370
rect 2974 430 2976 433
rect 3297 473 3299 500
rect 3318 473 3320 500
rect 3343 480 3345 500
rect 3161 455 3163 458
rect 3343 457 3345 460
rect 3297 430 3299 433
rect 3318 430 3320 433
rect 3073 407 3075 411
rect 3094 407 3096 411
rect 3115 407 3117 411
rect 2886 363 2888 366
rect 2907 363 2909 366
rect 2928 363 2930 366
rect 2949 363 2951 366
rect 2704 340 2706 343
rect 2725 340 2727 343
rect 2323 312 2325 319
rect 2318 308 2325 312
rect 2319 297 2321 308
rect 2331 300 2333 319
rect 2361 311 2363 319
rect 2405 311 2407 319
rect 2355 309 2363 311
rect 2399 309 2407 311
rect 2355 297 2357 309
rect 2363 297 2365 306
rect 2399 297 2401 309
rect 2407 297 2409 306
rect 2450 297 2452 319
rect 2319 284 2321 287
rect 2355 284 2357 287
rect 2363 284 2365 287
rect 2399 284 2401 287
rect 2407 284 2409 287
rect 2450 284 2452 287
rect 2898 282 2902 284
rect 2922 282 2949 284
rect 3109 282 3116 284
rect 3260 267 3262 271
rect 2898 261 2902 263
rect 2922 261 2949 263
rect 3109 261 3131 263
rect 2898 240 2902 242
rect 2922 240 2949 242
rect 3109 240 3144 242
rect 3373 266 3375 270
rect 3297 259 3299 266
rect 3330 252 3332 266
rect 3297 236 3299 239
rect 3330 229 3332 232
rect 2898 219 2902 221
rect 2922 219 2949 221
rect 3109 219 3155 221
rect 3260 207 3262 227
rect 3297 219 3299 222
rect 2906 194 2909 196
rect 2929 194 2949 196
rect 2989 194 3116 196
rect 3330 212 3332 215
rect 3260 184 3262 187
rect 3297 185 3299 199
rect 3373 206 3375 226
rect 3330 185 3332 192
rect 3373 183 3375 186
rect 3511 176 3513 179
rect 3519 176 3521 179
rect 3549 176 3551 179
rect 3593 176 3595 179
rect 3638 176 3640 179
rect 3511 144 3513 151
rect 3506 140 3513 144
rect 3507 129 3509 140
rect 3519 132 3521 151
rect 3549 143 3551 151
rect 3593 143 3595 151
rect 3543 141 3551 143
rect 3587 141 3595 143
rect 3543 129 3545 141
rect 3551 129 3553 138
rect 3587 129 3589 141
rect 3595 129 3597 138
rect 3638 129 3640 151
rect 3507 116 3509 119
rect 3543 116 3545 119
rect 3551 116 3553 119
rect 3587 116 3589 119
rect 3595 116 3597 119
rect 3638 116 3640 119
rect 2965 82 2967 85
rect 2973 82 2975 85
rect 3003 82 3005 85
rect 3047 82 3049 85
rect 3092 82 3094 85
rect 2965 50 2967 57
rect 2960 46 2967 50
rect 2961 35 2963 46
rect 2973 38 2975 57
rect 3003 49 3005 57
rect 3047 49 3049 57
rect 2997 47 3005 49
rect 3041 47 3049 49
rect 2997 35 2999 47
rect 3005 35 3007 44
rect 3041 35 3043 47
rect 3049 35 3051 44
rect 3092 35 3094 57
rect 2961 22 2963 25
rect 2997 22 2999 25
rect 3005 22 3007 25
rect 3041 22 3043 25
rect 3049 22 3051 25
rect 3092 22 3094 25
<< polycontact >>
rect 2247 1361 2251 1365
rect 2260 1353 2264 1357
rect 2271 1361 2275 1365
rect 2283 1353 2288 1358
rect 2298 1353 2302 1357
rect 2327 1353 2332 1358
rect 2379 1358 2383 1363
rect 2342 1353 2346 1357
rect 2718 1262 2724 1267
rect 2062 1254 2066 1258
rect 2025 1248 2029 1253
rect 2076 1253 2081 1258
rect 2106 1254 2110 1258
rect 2120 1253 2125 1258
rect 2133 1246 2137 1250
rect 2144 1254 2148 1258
rect 2157 1246 2161 1250
rect 2551 1244 2555 1249
rect 2584 1244 2588 1249
rect 2511 1188 2515 1193
rect 2253 1157 2257 1161
rect 2266 1149 2270 1153
rect 2277 1157 2281 1161
rect 2289 1149 2294 1154
rect 2304 1149 2308 1153
rect 2333 1149 2338 1154
rect 2385 1154 2389 1159
rect 2348 1149 2352 1153
rect 2624 1187 2628 1192
rect 2692 1183 2699 1189
rect 2741 1186 2745 1191
rect 2551 1158 2555 1163
rect 2584 1158 2588 1163
rect 2874 1207 2878 1212
rect 2907 1207 2911 1212
rect 2834 1151 2838 1156
rect 3113 1239 3117 1244
rect 3146 1239 3150 1244
rect 3073 1183 3077 1188
rect 2947 1150 2951 1155
rect 3186 1182 3190 1187
rect 3356 1169 3360 1173
rect 3113 1153 3117 1158
rect 3146 1153 3150 1158
rect 3369 1161 3373 1165
rect 3380 1169 3384 1173
rect 3392 1161 3397 1166
rect 3407 1161 3411 1165
rect 3436 1161 3441 1166
rect 3488 1166 3492 1171
rect 3451 1161 3455 1165
rect 2874 1121 2878 1126
rect 2907 1121 2911 1126
rect 2256 1028 2260 1032
rect 2269 1020 2273 1024
rect 2280 1028 2284 1032
rect 2292 1020 2297 1025
rect 2307 1020 2311 1024
rect 2336 1020 2341 1025
rect 2388 1025 2392 1030
rect 2351 1020 2355 1024
rect 3359 1033 3363 1037
rect 3372 1025 3376 1029
rect 3383 1033 3387 1037
rect 3395 1025 3400 1030
rect 3410 1025 3414 1029
rect 3439 1025 3444 1030
rect 3491 1030 3495 1035
rect 3454 1025 3458 1029
rect 3050 1007 3056 1012
rect 2934 1002 2940 1007
rect 2698 968 2704 973
rect 2531 950 2535 955
rect 2564 950 2568 955
rect 2491 894 2495 899
rect 2266 867 2270 871
rect 2279 859 2283 863
rect 2290 867 2294 871
rect 2302 859 2307 864
rect 2317 859 2321 863
rect 2346 859 2351 864
rect 2398 864 2402 869
rect 2361 859 2365 863
rect 2604 893 2608 898
rect 2908 923 2915 929
rect 2957 926 2961 931
rect 2672 889 2679 895
rect 2721 892 2725 897
rect 2531 864 2535 869
rect 2564 864 2568 869
rect 3024 891 3031 897
rect 3073 893 3077 898
rect 3317 851 3323 856
rect 3296 841 3302 846
rect 2937 792 2943 797
rect 3132 792 3138 797
rect 2916 779 2922 784
rect 2266 742 2270 746
rect 2279 734 2283 738
rect 2290 742 2294 746
rect 2302 734 2307 739
rect 2317 734 2321 738
rect 2346 734 2351 739
rect 2398 739 2402 744
rect 2361 734 2365 738
rect 2708 723 2714 728
rect 2541 705 2545 710
rect 2574 705 2578 710
rect 2501 649 2505 654
rect 2614 648 2618 653
rect 2890 700 2897 706
rect 2981 703 2985 708
rect 3106 713 3113 719
rect 3155 716 3159 721
rect 2682 644 2689 650
rect 2731 647 2735 652
rect 2541 619 2545 624
rect 2574 619 2578 624
rect 3270 681 3277 687
rect 3339 683 3343 688
rect 2266 576 2270 580
rect 2279 568 2283 572
rect 2290 576 2294 580
rect 2302 568 2307 573
rect 2317 568 2321 572
rect 2346 568 2351 573
rect 2398 573 2402 578
rect 2361 568 2365 572
rect 2947 570 2953 575
rect 3113 570 3119 575
rect 2926 559 2932 564
rect 2905 532 2911 537
rect 3092 559 3098 564
rect 3316 559 3322 564
rect 2723 469 2729 474
rect 3066 478 3073 484
rect 2266 451 2270 455
rect 2279 443 2283 447
rect 2290 451 2294 455
rect 2302 443 2307 448
rect 2317 443 2321 447
rect 2346 443 2351 448
rect 2398 448 2402 453
rect 2361 443 2365 447
rect 2556 451 2560 456
rect 2589 451 2593 456
rect 2516 395 2520 400
rect 2879 453 2886 459
rect 2629 394 2633 399
rect 2970 456 2974 461
rect 3157 481 3161 486
rect 3290 480 3297 486
rect 2697 390 2704 396
rect 2746 393 2750 398
rect 2556 365 2560 370
rect 2589 365 2593 370
rect 3339 483 3343 488
rect 2314 308 2318 312
rect 2327 300 2331 304
rect 2338 308 2342 312
rect 2350 300 2355 305
rect 2365 300 2369 304
rect 2394 300 2399 305
rect 2446 305 2450 310
rect 2409 300 2413 304
rect 2929 284 2935 291
rect 3131 259 3136 265
rect 3144 238 3149 244
rect 3296 266 3300 271
rect 3329 266 3333 271
rect 3155 217 3160 223
rect 3256 210 3260 215
rect 2932 196 2937 200
rect 3369 209 3373 214
rect 3296 180 3300 185
rect 3329 180 3333 185
rect 3502 140 3506 144
rect 3515 132 3519 136
rect 3526 140 3530 144
rect 3538 132 3543 137
rect 3553 132 3557 136
rect 3582 132 3587 137
rect 3634 137 3638 142
rect 3597 132 3601 136
rect 2956 46 2960 50
rect 2969 38 2973 42
rect 2980 46 2984 50
rect 2992 38 2997 43
rect 3007 38 3011 42
rect 3036 38 3041 43
rect 3088 43 3092 48
rect 3051 38 3055 42
<< metal1 >>
rect 2244 1403 2398 1408
rect 2251 1397 2255 1403
rect 2289 1397 2293 1403
rect 2333 1397 2337 1403
rect 2378 1397 2382 1403
rect 2301 1372 2314 1397
rect 2345 1372 2358 1397
rect 2240 1361 2247 1365
rect 2251 1353 2260 1357
rect 2267 1350 2271 1372
rect 2275 1361 2276 1365
rect 2311 1363 2314 1372
rect 2355 1363 2358 1372
rect 2311 1358 2323 1363
rect 2355 1358 2379 1363
rect 2386 1362 2390 1372
rect 2275 1356 2283 1358
rect 2280 1353 2283 1356
rect 2302 1353 2303 1357
rect 2311 1350 2314 1358
rect 2319 1353 2327 1358
rect 2346 1353 2347 1357
rect 2355 1350 2358 1358
rect 2386 1357 2403 1362
rect 2386 1350 2390 1357
rect 2259 1340 2271 1350
rect 2303 1340 2314 1350
rect 2347 1340 2358 1350
rect 2247 1335 2251 1340
rect 2283 1335 2287 1340
rect 2327 1335 2331 1340
rect 2378 1335 2382 1340
rect 2246 1331 2390 1335
rect 2399 1302 2403 1357
rect 2005 1254 2009 1300
rect 2399 1297 2708 1302
rect 2495 1281 2757 1286
rect 2018 1276 2162 1280
rect 2026 1271 2030 1276
rect 2077 1271 2081 1276
rect 2121 1271 2125 1276
rect 2157 1271 2161 1276
rect 2050 1261 2061 1271
rect 2094 1261 2105 1271
rect 2137 1261 2149 1271
rect 2018 1254 2022 1261
rect 2005 1249 2022 1254
rect 2050 1253 2053 1261
rect 2061 1254 2062 1258
rect 2081 1253 2089 1258
rect 2094 1253 2097 1261
rect 2105 1254 2106 1258
rect 2125 1255 2128 1258
rect 2125 1253 2133 1255
rect 2018 1239 2022 1249
rect 2029 1248 2053 1253
rect 2085 1248 2097 1253
rect 2050 1239 2053 1248
rect 2094 1239 2097 1248
rect 2132 1246 2133 1250
rect 2137 1239 2141 1261
rect 2148 1254 2157 1258
rect 2161 1246 2171 1250
rect 2050 1214 2063 1239
rect 2094 1214 2107 1239
rect 2168 1230 2171 1246
rect 2510 1245 2514 1281
rect 2168 1226 2475 1230
rect 2026 1208 2030 1214
rect 2071 1208 2075 1214
rect 2115 1208 2119 1214
rect 2153 1208 2157 1214
rect 2010 1203 2164 1208
rect 2250 1199 2404 1204
rect 2257 1193 2261 1199
rect 2295 1193 2299 1199
rect 2339 1193 2343 1199
rect 2384 1193 2388 1199
rect 2307 1168 2320 1193
rect 2351 1168 2364 1193
rect 2246 1157 2253 1161
rect 2257 1149 2266 1153
rect 2273 1146 2277 1168
rect 2281 1157 2282 1161
rect 2317 1159 2320 1168
rect 2361 1159 2364 1168
rect 2317 1154 2329 1159
rect 2361 1154 2385 1159
rect 2392 1158 2396 1168
rect 2281 1152 2289 1154
rect 2286 1149 2289 1152
rect 2308 1149 2309 1153
rect 2317 1146 2320 1154
rect 2325 1149 2333 1154
rect 2352 1149 2353 1153
rect 2361 1146 2364 1154
rect 2392 1153 2408 1158
rect 2392 1146 2396 1153
rect 2265 1136 2277 1146
rect 2309 1136 2320 1146
rect 2353 1136 2364 1146
rect 2253 1131 2257 1136
rect 2289 1131 2293 1136
rect 2333 1131 2337 1136
rect 2384 1131 2388 1136
rect 2252 1127 2396 1131
rect 2405 1103 2408 1153
rect 2470 1150 2475 1226
rect 2535 1213 2540 1268
rect 2551 1249 2555 1256
rect 2584 1249 2588 1256
rect 2623 1244 2627 1281
rect 2670 1262 2708 1267
rect 2714 1262 2718 1267
rect 2724 1262 2726 1267
rect 2670 1261 2681 1262
rect 2643 1256 2681 1261
rect 2751 1256 2757 1281
rect 3044 1276 3277 1281
rect 2688 1248 2759 1256
rect 2777 1254 3048 1259
rect 2547 1213 2551 1217
rect 2535 1209 2551 1213
rect 2501 1188 2511 1193
rect 2518 1192 2522 1205
rect 2547 1197 2551 1209
rect 2518 1187 2531 1192
rect 2518 1185 2522 1187
rect 2555 1212 2559 1217
rect 2555 1208 2573 1212
rect 2555 1197 2559 1208
rect 2568 1198 2573 1208
rect 2580 1198 2584 1210
rect 2568 1194 2584 1198
rect 2569 1193 2584 1194
rect 2510 1126 2514 1165
rect 2551 1145 2555 1158
rect 2569 1135 2574 1193
rect 2580 1190 2584 1193
rect 2588 1197 2592 1210
rect 2588 1193 2609 1197
rect 2588 1190 2592 1193
rect 2603 1192 2609 1193
rect 2603 1187 2613 1192
rect 2619 1187 2624 1192
rect 2631 1191 2635 1204
rect 2694 1243 2698 1248
rect 2723 1243 2727 1248
rect 2740 1243 2744 1248
rect 2631 1186 2648 1191
rect 2631 1184 2635 1186
rect 2673 1183 2692 1189
rect 2707 1184 2712 1203
rect 2733 1186 2741 1191
rect 2748 1190 2752 1203
rect 2777 1190 2781 1254
rect 2805 1244 3038 1249
rect 2733 1184 2737 1186
rect 2584 1145 2588 1158
rect 2623 1126 2627 1164
rect 2673 1146 2681 1183
rect 2707 1180 2737 1184
rect 2748 1185 2781 1190
rect 2748 1183 2752 1185
rect 2723 1176 2727 1180
rect 2740 1146 2744 1163
rect 2733 1143 2744 1146
rect 2694 1126 2698 1136
rect 2733 1126 2739 1143
rect 2495 1118 2750 1126
rect 2405 1094 2673 1103
rect 2405 1093 2408 1094
rect 2253 1070 2407 1075
rect 2260 1064 2264 1070
rect 2298 1064 2302 1070
rect 2342 1064 2346 1070
rect 2387 1064 2391 1070
rect 2310 1039 2323 1064
rect 2354 1039 2367 1064
rect 2249 1028 2256 1032
rect 2260 1020 2269 1024
rect 2276 1017 2280 1039
rect 2284 1028 2285 1032
rect 2320 1030 2323 1039
rect 2364 1030 2367 1039
rect 2395 1030 2399 1039
rect 2320 1025 2332 1030
rect 2364 1025 2388 1030
rect 2284 1023 2292 1025
rect 2289 1020 2292 1023
rect 2311 1020 2312 1024
rect 2320 1017 2323 1025
rect 2328 1020 2336 1025
rect 2355 1020 2356 1024
rect 2364 1017 2367 1025
rect 2395 1024 2681 1030
rect 2395 1017 2399 1024
rect 2268 1007 2280 1017
rect 2312 1007 2323 1017
rect 2356 1007 2367 1017
rect 2678 1008 2681 1024
rect 2256 1002 2260 1007
rect 2292 1002 2296 1007
rect 2336 1002 2340 1007
rect 2387 1002 2391 1007
rect 2678 1003 2688 1008
rect 2777 1007 2781 1185
rect 2833 1208 2837 1244
rect 2858 1176 2863 1231
rect 2874 1212 2878 1219
rect 2907 1212 2911 1219
rect 2946 1207 2950 1244
rect 3044 1230 3048 1254
rect 2993 1224 3048 1230
rect 2966 1219 3048 1224
rect 3072 1240 3076 1276
rect 2870 1176 2874 1180
rect 2858 1172 2874 1176
rect 2824 1151 2834 1156
rect 2841 1155 2845 1168
rect 2870 1160 2874 1172
rect 2841 1150 2854 1155
rect 2841 1148 2845 1150
rect 2878 1175 2882 1180
rect 2878 1171 2895 1175
rect 2878 1160 2882 1171
rect 2891 1161 2895 1171
rect 2903 1161 2907 1173
rect 2891 1156 2907 1161
rect 2833 1089 2837 1128
rect 2874 1108 2878 1121
rect 2891 1099 2897 1156
rect 2903 1153 2907 1156
rect 2911 1160 2915 1173
rect 3097 1208 3102 1263
rect 3113 1244 3117 1251
rect 3146 1244 3150 1251
rect 3185 1239 3189 1276
rect 3232 1256 3283 1262
rect 3205 1251 3283 1256
rect 3109 1208 3113 1212
rect 3097 1204 3113 1208
rect 3063 1183 3073 1188
rect 3080 1187 3084 1200
rect 3109 1192 3113 1204
rect 3080 1182 3093 1187
rect 3080 1180 3084 1182
rect 2911 1156 2932 1160
rect 2911 1153 2915 1156
rect 2926 1155 2932 1156
rect 2926 1150 2936 1155
rect 2942 1150 2947 1155
rect 2954 1154 2958 1167
rect 3117 1207 3121 1212
rect 3117 1203 3134 1207
rect 3117 1192 3121 1203
rect 3130 1193 3134 1203
rect 3142 1193 3146 1205
rect 3130 1188 3146 1193
rect 2954 1149 2971 1154
rect 2954 1147 2958 1149
rect 2996 1146 3036 1152
rect 2907 1108 2911 1121
rect 2946 1089 2950 1127
rect 2996 1109 3004 1146
rect 2805 1081 3014 1089
rect 3028 1049 3036 1146
rect 3072 1121 3076 1160
rect 3113 1140 3117 1153
rect 3130 1131 3136 1188
rect 3142 1185 3146 1188
rect 3150 1192 3154 1205
rect 3353 1211 3507 1216
rect 3150 1188 3171 1192
rect 3150 1185 3154 1188
rect 3165 1187 3171 1188
rect 3165 1182 3175 1187
rect 3181 1182 3186 1187
rect 3193 1186 3197 1199
rect 3360 1205 3364 1211
rect 3398 1205 3402 1211
rect 3442 1205 3446 1211
rect 3487 1205 3491 1211
rect 3193 1181 3210 1186
rect 3193 1179 3197 1181
rect 3235 1178 3272 1184
rect 3410 1180 3423 1205
rect 3454 1180 3467 1205
rect 3146 1140 3150 1153
rect 3185 1121 3189 1159
rect 3235 1141 3243 1178
rect 3044 1113 3253 1121
rect 3268 1107 3272 1178
rect 3288 1169 3356 1173
rect 3360 1161 3369 1165
rect 3376 1158 3380 1180
rect 3384 1169 3385 1173
rect 3420 1171 3423 1180
rect 3464 1171 3467 1180
rect 3420 1166 3432 1171
rect 3464 1166 3488 1171
rect 3495 1170 3499 1180
rect 3384 1164 3392 1166
rect 3389 1161 3392 1164
rect 3411 1161 3412 1165
rect 3420 1158 3423 1166
rect 3428 1161 3436 1166
rect 3455 1161 3456 1165
rect 3464 1158 3467 1166
rect 3495 1165 3512 1170
rect 3495 1158 3499 1165
rect 3368 1148 3380 1158
rect 3412 1148 3423 1158
rect 3456 1148 3467 1158
rect 3356 1143 3360 1148
rect 3392 1143 3396 1148
rect 3436 1143 3440 1148
rect 3487 1143 3491 1148
rect 3355 1139 3499 1143
rect 3508 1122 3512 1165
rect 2804 1043 3036 1049
rect 2906 1031 3116 1034
rect 2906 1026 3098 1031
rect 3104 1026 3116 1031
rect 2906 1024 3091 1026
rect 2906 1023 2975 1024
rect 2777 1002 2865 1007
rect 2870 1002 2934 1007
rect 2255 998 2399 1002
rect 2967 996 2975 1023
rect 2987 1007 3050 1012
rect 3083 1001 3091 1024
rect 2475 987 2737 992
rect 2903 988 2975 996
rect 3019 993 3091 1001
rect 3026 990 3030 993
rect 2490 951 2494 987
rect 2263 909 2417 914
rect 2515 919 2520 974
rect 2531 955 2535 962
rect 2564 955 2568 962
rect 2603 950 2607 987
rect 2650 968 2688 973
rect 2694 968 2698 973
rect 2704 968 2706 973
rect 2650 967 2661 968
rect 2623 962 2661 967
rect 2731 962 2737 987
rect 2910 983 2914 988
rect 2939 983 2943 988
rect 2668 954 2739 962
rect 2527 919 2531 923
rect 2515 915 2531 919
rect 2270 903 2274 909
rect 2308 903 2312 909
rect 2352 903 2356 909
rect 2397 903 2401 909
rect 2320 878 2333 903
rect 2364 878 2377 903
rect 2481 894 2491 899
rect 2498 898 2502 911
rect 2527 903 2531 915
rect 2498 893 2511 898
rect 2498 891 2502 893
rect 2259 867 2266 871
rect 2270 859 2279 863
rect 2286 856 2290 878
rect 2294 867 2295 871
rect 2330 869 2333 878
rect 2374 869 2377 878
rect 2330 864 2342 869
rect 2374 864 2398 869
rect 2405 868 2409 878
rect 2535 918 2539 923
rect 2535 914 2553 918
rect 2535 903 2539 914
rect 2548 904 2553 914
rect 2560 904 2564 916
rect 2548 900 2564 904
rect 2549 899 2564 900
rect 2294 862 2302 864
rect 2299 859 2302 862
rect 2321 859 2322 863
rect 2330 856 2333 864
rect 2338 859 2346 864
rect 2365 859 2366 863
rect 2374 856 2377 864
rect 2405 863 2423 868
rect 2405 856 2409 863
rect 2278 846 2290 856
rect 2322 846 2333 856
rect 2366 846 2377 856
rect 2266 841 2270 846
rect 2302 841 2306 846
rect 2346 841 2350 846
rect 2397 841 2401 846
rect 2265 837 2409 841
rect 2418 809 2423 863
rect 2490 832 2494 871
rect 2531 851 2535 864
rect 2549 841 2554 899
rect 2560 896 2564 899
rect 2568 903 2572 916
rect 2568 899 2589 903
rect 2568 896 2572 899
rect 2583 898 2589 899
rect 2583 893 2593 898
rect 2599 893 2604 898
rect 2611 897 2615 910
rect 2674 949 2678 954
rect 2703 949 2707 954
rect 2720 949 2724 954
rect 2956 983 2960 988
rect 2792 923 2874 929
rect 2879 923 2908 929
rect 2923 924 2928 943
rect 2949 926 2957 931
rect 2964 930 2968 943
rect 2949 924 2953 926
rect 2923 920 2953 924
rect 2964 925 2982 930
rect 2964 923 2968 925
rect 2939 916 2943 920
rect 2611 892 2628 897
rect 2611 890 2615 892
rect 2653 889 2672 895
rect 2687 890 2692 909
rect 2713 892 2721 897
rect 2728 896 2732 909
rect 2713 890 2717 892
rect 2564 851 2568 864
rect 2603 832 2607 870
rect 2653 852 2661 889
rect 2687 886 2717 890
rect 2728 891 2761 896
rect 2728 889 2732 891
rect 2703 882 2707 886
rect 2720 852 2724 869
rect 2713 849 2724 852
rect 2674 832 2678 842
rect 2713 832 2719 849
rect 2756 845 2761 891
rect 3038 910 3047 990
rect 3072 950 3076 993
rect 2956 886 2960 903
rect 3055 898 3059 910
rect 2982 891 3024 897
rect 3039 893 3073 898
rect 3080 897 3084 910
rect 3268 897 3272 1102
rect 3356 1075 3510 1080
rect 3363 1069 3367 1075
rect 3401 1069 3405 1075
rect 3445 1069 3449 1075
rect 3490 1069 3494 1075
rect 3291 1037 3296 1064
rect 3413 1044 3426 1069
rect 3457 1044 3470 1069
rect 3291 1033 3359 1037
rect 3363 1025 3372 1029
rect 3379 1022 3383 1044
rect 3387 1033 3388 1037
rect 3423 1035 3426 1044
rect 3467 1035 3470 1044
rect 3423 1030 3435 1035
rect 3467 1030 3491 1035
rect 3498 1034 3502 1044
rect 3387 1028 3395 1030
rect 3392 1025 3395 1028
rect 3414 1025 3415 1029
rect 3423 1022 3426 1030
rect 3431 1025 3439 1030
rect 3458 1025 3459 1029
rect 3467 1022 3470 1030
rect 3498 1029 3515 1034
rect 3498 1022 3502 1029
rect 3371 1012 3383 1022
rect 3415 1012 3426 1022
rect 3459 1012 3470 1022
rect 3359 1007 3363 1012
rect 3395 1007 3399 1012
rect 3439 1007 3443 1012
rect 3490 1007 3494 1012
rect 3358 1003 3502 1007
rect 3511 986 3515 1029
rect 3039 888 3044 893
rect 3080 892 3306 897
rect 3080 890 3084 892
rect 2949 883 2960 886
rect 2910 866 2914 876
rect 2949 866 2955 883
rect 3038 868 3047 888
rect 2900 864 2961 866
rect 3026 864 3030 868
rect 3055 864 3059 868
rect 3072 864 3076 870
rect 2900 858 3036 864
rect 3043 858 3109 864
rect 3215 860 3383 868
rect 3390 860 3391 868
rect 3238 851 3317 856
rect 2756 839 3076 845
rect 2475 824 2730 832
rect 3054 814 3098 819
rect 3104 814 3225 819
rect 3054 811 3225 814
rect 2418 800 2653 809
rect 2887 803 3059 811
rect 2845 792 2874 797
rect 2879 792 2937 797
rect 2943 792 3132 797
rect 2263 784 2417 789
rect 3165 786 3173 811
rect 3238 805 3244 851
rect 2270 778 2274 784
rect 2308 778 2312 784
rect 2352 778 2356 784
rect 2397 778 2401 784
rect 2791 779 2853 784
rect 2858 779 2916 784
rect 3101 778 3173 786
rect 3189 801 3244 805
rect 3252 841 3296 846
rect 2320 753 2333 778
rect 2364 753 2377 778
rect 3108 773 3112 778
rect 3137 773 3141 778
rect 2885 765 2999 773
rect 2259 742 2266 746
rect 2270 734 2279 738
rect 2286 731 2290 753
rect 2294 742 2295 746
rect 2330 744 2333 753
rect 2374 744 2377 753
rect 2330 739 2342 744
rect 2374 739 2398 744
rect 2405 743 2409 753
rect 2424 758 2698 763
rect 2892 760 2896 765
rect 2928 760 2932 765
rect 2980 760 2984 765
rect 2424 743 2428 758
rect 2294 737 2302 739
rect 2299 734 2302 737
rect 2321 734 2322 738
rect 2330 731 2333 739
rect 2338 734 2346 739
rect 2365 734 2366 738
rect 2374 731 2377 739
rect 2405 738 2428 743
rect 2485 742 2747 747
rect 2405 731 2409 738
rect 2278 721 2290 731
rect 2322 721 2333 731
rect 2366 721 2377 731
rect 2266 716 2270 721
rect 2302 716 2306 721
rect 2346 716 2350 721
rect 2397 716 2401 721
rect 2265 712 2409 716
rect 2500 706 2504 742
rect 2525 674 2530 729
rect 2541 710 2545 717
rect 2574 710 2578 717
rect 2613 705 2617 742
rect 2660 723 2698 728
rect 2704 723 2708 728
rect 2714 723 2716 728
rect 2660 722 2671 723
rect 2633 717 2671 722
rect 2741 717 2747 742
rect 3154 773 3158 778
rect 2678 709 2749 717
rect 2537 674 2541 678
rect 2525 670 2541 674
rect 2491 649 2501 654
rect 2508 653 2512 666
rect 2537 658 2541 670
rect 2508 648 2521 653
rect 2508 646 2512 648
rect 2545 673 2549 678
rect 2545 669 2563 673
rect 2545 658 2549 669
rect 2558 659 2563 669
rect 2570 659 2574 671
rect 2558 655 2574 659
rect 2559 654 2574 655
rect 2263 618 2417 623
rect 2270 612 2274 618
rect 2308 612 2312 618
rect 2352 612 2356 618
rect 2397 612 2401 618
rect 2320 587 2333 612
rect 2364 587 2377 612
rect 2500 587 2504 626
rect 2541 606 2545 619
rect 2559 596 2564 654
rect 2570 651 2574 654
rect 2578 658 2582 671
rect 2578 654 2599 658
rect 2578 651 2582 654
rect 2593 653 2599 654
rect 2593 648 2603 653
rect 2609 648 2614 653
rect 2621 652 2625 665
rect 2684 704 2688 709
rect 2713 704 2717 709
rect 2730 704 2734 709
rect 2870 700 2890 706
rect 2905 701 2909 720
rect 2942 701 2946 720
rect 2973 703 2981 708
rect 2988 707 2992 720
rect 3029 713 3076 719
rect 3083 713 3106 719
rect 3121 714 3126 733
rect 3147 716 3155 721
rect 3162 720 3166 733
rect 3189 720 3193 801
rect 3147 714 3151 716
rect 3121 710 3151 714
rect 3162 715 3193 720
rect 3162 713 3166 715
rect 2973 701 2977 703
rect 2905 697 2977 701
rect 2988 702 3082 707
rect 3137 706 3141 710
rect 2988 700 2992 702
rect 2942 693 2946 697
rect 2621 647 2638 652
rect 2621 645 2625 647
rect 2663 644 2682 650
rect 2697 645 2702 664
rect 2723 647 2731 652
rect 2738 651 2742 664
rect 2723 645 2727 647
rect 2574 606 2578 619
rect 2613 587 2617 625
rect 2663 607 2671 644
rect 2697 641 2727 645
rect 2738 646 2771 651
rect 2738 644 2742 646
rect 2713 637 2717 641
rect 2730 607 2734 624
rect 2723 604 2734 607
rect 2765 607 2771 646
rect 2904 633 2913 693
rect 2925 633 2934 693
rect 2980 653 2984 680
rect 3252 708 3258 841
rect 3349 835 3357 860
rect 3265 827 3357 835
rect 3272 819 3276 827
rect 3284 699 3293 819
rect 3305 699 3314 819
rect 3338 740 3342 827
rect 3154 676 3158 693
rect 3322 688 3326 699
rect 3242 681 3270 687
rect 3285 683 3339 688
rect 3346 687 3350 700
rect 3285 678 3290 683
rect 3322 678 3326 683
rect 3346 682 3405 687
rect 3346 680 3350 682
rect 3147 673 3158 676
rect 3108 653 3112 666
rect 3147 653 3151 673
rect 3284 658 3293 678
rect 3305 658 3314 678
rect 3272 653 3276 658
rect 3307 653 3311 658
rect 3338 653 3342 660
rect 2980 648 3036 653
rect 3043 648 3217 653
rect 3227 648 3391 653
rect 2892 622 2896 633
rect 2980 622 2984 648
rect 2883 614 2984 622
rect 2684 587 2688 597
rect 2723 587 2729 604
rect 2765 602 3236 607
rect 2259 576 2266 580
rect 2270 568 2279 572
rect 2286 565 2290 587
rect 2294 576 2295 580
rect 2330 578 2333 587
rect 2374 578 2377 587
rect 2330 573 2342 578
rect 2374 573 2398 578
rect 2405 577 2409 587
rect 2485 579 2740 587
rect 2878 581 3197 589
rect 3206 586 3249 589
rect 3206 581 3383 586
rect 3235 578 3383 581
rect 3390 578 3391 586
rect 2294 571 2302 573
rect 2299 568 2302 571
rect 2321 568 2322 572
rect 2330 565 2333 573
rect 2338 568 2346 573
rect 2365 568 2366 572
rect 2374 565 2377 573
rect 2405 572 2418 577
rect 2405 565 2409 572
rect 2414 569 2418 572
rect 2858 570 2947 575
rect 2953 570 3113 575
rect 2414 565 2655 569
rect 2278 555 2290 565
rect 2322 555 2333 565
rect 2366 555 2377 565
rect 2649 564 2655 565
rect 2649 555 2663 564
rect 2803 559 2926 564
rect 2932 559 3092 564
rect 3098 559 3316 564
rect 2266 550 2270 555
rect 2302 550 2306 555
rect 2346 550 2350 555
rect 2397 550 2401 555
rect 3349 553 3357 578
rect 2265 546 2409 550
rect 3061 543 3175 551
rect 3285 545 3357 553
rect 3068 538 3072 543
rect 3104 538 3108 543
rect 3156 538 3160 543
rect 3292 540 3296 545
rect 3321 540 3325 545
rect 2870 532 2905 537
rect 2874 518 2988 526
rect 2881 513 2885 518
rect 2916 513 2920 518
rect 2952 513 2956 518
rect 2430 504 2713 509
rect 2263 493 2417 498
rect 2270 487 2274 493
rect 2308 487 2312 493
rect 2352 487 2356 493
rect 2397 487 2401 493
rect 2320 462 2333 487
rect 2364 462 2377 487
rect 2259 451 2266 455
rect 2270 443 2279 447
rect 2286 440 2290 462
rect 2294 451 2295 455
rect 2330 453 2333 462
rect 2374 453 2377 462
rect 2330 448 2342 453
rect 2374 448 2398 453
rect 2405 452 2409 462
rect 2430 452 2434 504
rect 2500 488 2762 493
rect 2294 446 2302 448
rect 2299 443 2302 446
rect 2321 443 2322 447
rect 2330 440 2333 448
rect 2338 443 2346 448
rect 2365 443 2366 447
rect 2374 440 2377 448
rect 2405 447 2434 452
rect 2515 452 2519 488
rect 2405 440 2409 447
rect 2278 430 2290 440
rect 2322 430 2333 440
rect 2366 430 2377 440
rect 2266 425 2270 430
rect 2302 425 2306 430
rect 2346 425 2350 430
rect 2397 425 2401 430
rect 2265 421 2409 425
rect 2540 420 2545 475
rect 2556 456 2560 463
rect 2589 456 2593 463
rect 2628 451 2632 488
rect 2675 469 2713 474
rect 2719 469 2723 474
rect 2729 469 2731 474
rect 2675 468 2686 469
rect 2648 463 2686 468
rect 2756 463 2762 488
rect 2969 513 2973 518
rect 3338 540 3342 545
rect 3029 478 3066 484
rect 3081 479 3085 498
rect 3118 479 3122 498
rect 3149 481 3157 486
rect 3164 485 3168 498
rect 3149 479 3153 481
rect 3081 475 3153 479
rect 3164 480 3176 485
rect 3242 480 3290 486
rect 3305 481 3310 500
rect 3331 483 3339 488
rect 3346 487 3350 500
rect 3331 481 3335 483
rect 3164 478 3168 480
rect 2693 455 2764 463
rect 2552 420 2556 424
rect 2540 416 2556 420
rect 2506 395 2516 400
rect 2523 399 2527 412
rect 2552 404 2556 416
rect 2523 394 2536 399
rect 2523 392 2527 394
rect 2560 419 2564 424
rect 2560 415 2578 419
rect 2560 404 2564 415
rect 2573 405 2578 415
rect 2585 405 2589 417
rect 2573 401 2589 405
rect 2574 400 2589 401
rect 2311 350 2465 355
rect 2318 344 2322 350
rect 2356 344 2360 350
rect 2400 344 2404 350
rect 2445 344 2449 350
rect 2368 319 2381 344
rect 2412 319 2425 344
rect 2515 333 2519 372
rect 2556 352 2560 365
rect 2574 342 2579 400
rect 2585 397 2589 400
rect 2593 404 2597 417
rect 2593 400 2614 404
rect 2593 397 2597 400
rect 2608 399 2614 400
rect 2608 394 2618 399
rect 2624 394 2629 399
rect 2636 398 2640 411
rect 2699 450 2703 455
rect 2728 450 2732 455
rect 2745 450 2749 455
rect 2845 453 2879 459
rect 2894 454 2898 473
rect 2937 454 2941 473
rect 2962 456 2970 461
rect 2977 460 2981 473
rect 3118 471 3122 475
rect 2962 454 2966 456
rect 2894 450 2966 454
rect 2977 455 3013 460
rect 2977 453 2981 455
rect 2952 446 2956 450
rect 2636 393 2653 398
rect 2636 391 2640 393
rect 2678 390 2697 396
rect 2712 391 2717 410
rect 2738 393 2746 398
rect 2753 397 2757 410
rect 2738 391 2742 393
rect 2589 352 2593 365
rect 2628 333 2632 371
rect 2678 353 2686 390
rect 2712 387 2742 391
rect 2753 392 2786 397
rect 2753 390 2757 392
rect 2728 383 2732 387
rect 2745 353 2749 370
rect 2738 350 2749 353
rect 2699 333 2703 343
rect 2738 333 2744 350
rect 2781 333 2786 392
rect 2893 366 2902 446
rect 2914 366 2923 446
rect 2935 366 2944 446
rect 2969 378 2973 433
rect 3080 411 3089 471
rect 3101 411 3110 471
rect 3305 477 3335 481
rect 3346 482 3381 487
rect 3346 480 3350 482
rect 3321 473 3325 477
rect 3156 423 3160 458
rect 3338 443 3342 460
rect 3331 440 3342 443
rect 3292 423 3296 433
rect 3331 423 3337 440
rect 3156 415 3218 423
rect 3227 415 3356 423
rect 3068 378 3072 411
rect 3156 378 3160 415
rect 2969 370 3160 378
rect 2881 353 2885 366
rect 2969 353 2973 370
rect 2823 345 2973 353
rect 2500 325 2755 333
rect 2781 328 2873 333
rect 2307 308 2314 312
rect 2318 300 2327 304
rect 2334 297 2338 319
rect 2342 308 2343 312
rect 2378 310 2381 319
rect 2422 310 2425 319
rect 2378 305 2390 310
rect 2422 305 2446 310
rect 2453 309 2457 319
rect 2670 309 2678 310
rect 2342 303 2350 305
rect 2347 300 2350 303
rect 2369 300 2370 304
rect 2378 297 2381 305
rect 2386 300 2394 305
rect 2413 300 2414 304
rect 2422 297 2425 305
rect 2453 302 2678 309
rect 2453 297 2457 302
rect 2670 301 2678 302
rect 2326 287 2338 297
rect 2370 287 2381 297
rect 2414 287 2425 297
rect 2883 289 2891 345
rect 3378 333 3381 482
rect 2929 291 2935 333
rect 2314 282 2318 287
rect 2350 282 2354 287
rect 2394 282 2398 287
rect 2445 282 2449 287
rect 2883 285 2902 289
rect 2313 278 2457 282
rect 2883 254 2891 285
rect 3117 289 3125 296
rect 3109 285 3125 289
rect 2902 276 2922 277
rect 2902 271 2930 276
rect 2902 268 2922 271
rect 2902 254 2922 256
rect 2883 250 2922 254
rect 2883 218 2891 250
rect 2902 247 2922 250
rect 2902 232 2922 235
rect 2926 232 2930 271
rect 2949 268 3109 277
rect 2949 247 3109 256
rect 2902 228 2930 232
rect 2902 226 2922 228
rect 2926 218 2930 228
rect 2949 226 3109 235
rect 2883 214 2902 218
rect 2926 214 2949 218
rect 2883 201 2891 214
rect 2926 208 2930 214
rect 2926 204 2937 208
rect 2883 197 2909 201
rect 2932 200 2937 204
rect 3117 201 3125 285
rect 3131 265 3136 327
rect 3144 244 3149 327
rect 3155 327 3381 333
rect 3401 328 3405 682
rect 3155 223 3160 327
rect 3401 323 3471 328
rect 3227 303 3460 308
rect 2883 157 2891 197
rect 2989 197 3125 201
rect 2929 189 2949 193
rect 3117 190 3125 197
rect 3180 190 3188 303
rect 3255 267 3259 303
rect 3280 235 3285 290
rect 3296 271 3300 278
rect 3329 271 3333 278
rect 3368 266 3372 303
rect 3466 289 3471 323
rect 3415 283 3471 289
rect 3388 278 3471 283
rect 3292 235 3296 239
rect 3280 231 3296 235
rect 3246 210 3256 215
rect 3263 214 3267 227
rect 3292 219 3296 231
rect 3263 209 3276 214
rect 3263 207 3267 209
rect 2931 50 2936 189
rect 3117 179 3188 190
rect 3300 234 3304 239
rect 3300 230 3317 234
rect 3300 219 3304 230
rect 3313 220 3317 230
rect 3325 220 3329 232
rect 3313 215 3329 220
rect 3255 148 3259 187
rect 3296 167 3300 180
rect 3313 158 3319 215
rect 3325 212 3329 215
rect 3333 219 3337 232
rect 3333 215 3354 219
rect 3333 212 3337 215
rect 3348 214 3354 215
rect 3348 209 3358 214
rect 3364 209 3369 214
rect 3376 213 3380 226
rect 3376 208 3393 213
rect 3376 206 3380 208
rect 3418 205 3450 211
rect 3329 167 3333 180
rect 3368 148 3372 186
rect 3418 168 3426 205
rect 3499 182 3653 187
rect 3506 176 3510 182
rect 3544 176 3548 182
rect 3588 176 3592 182
rect 3633 176 3637 182
rect 3556 151 3569 176
rect 3600 151 3613 176
rect 3227 140 3436 148
rect 3474 140 3502 144
rect 3506 132 3515 136
rect 3522 129 3526 151
rect 3530 140 3531 144
rect 3566 142 3569 151
rect 3610 142 3613 151
rect 3566 137 3578 142
rect 3610 137 3634 142
rect 3641 141 3645 151
rect 3530 135 3538 137
rect 3535 132 3538 135
rect 3557 132 3558 136
rect 3566 129 3569 137
rect 3574 132 3582 137
rect 3601 132 3602 136
rect 3610 129 3613 137
rect 3641 136 3658 141
rect 3641 129 3645 136
rect 3514 119 3526 129
rect 3558 119 3569 129
rect 3602 119 3613 129
rect 3502 114 3506 119
rect 3538 114 3542 119
rect 3582 114 3586 119
rect 3633 114 3637 119
rect 3501 110 3645 114
rect 3654 94 3658 136
rect 2953 88 3107 93
rect 2960 82 2964 88
rect 2998 82 3002 88
rect 3042 82 3046 88
rect 3087 82 3091 88
rect 3010 57 3023 82
rect 3054 57 3067 82
rect 2931 46 2956 50
rect 2960 38 2969 42
rect 2976 35 2980 57
rect 2984 46 2985 50
rect 3020 48 3023 57
rect 3064 48 3067 57
rect 3020 43 3032 48
rect 3064 43 3088 48
rect 3095 47 3099 57
rect 2984 41 2992 43
rect 2989 38 2992 41
rect 3011 38 3012 42
rect 3020 35 3023 43
rect 3028 38 3036 43
rect 3055 38 3056 42
rect 3064 35 3067 43
rect 3095 42 3112 47
rect 3095 35 3099 42
rect 2968 25 2980 35
rect 3012 25 3023 35
rect 3056 25 3067 35
rect 2956 20 2960 25
rect 2992 20 2996 25
rect 3036 20 3040 25
rect 3087 20 3091 25
rect 2955 16 3099 20
rect 3108 -1 3112 42
<< m2contact >>
rect 2246 1353 2251 1358
rect 2276 1361 2281 1366
rect 2275 1351 2280 1356
rect 2303 1353 2308 1358
rect 2347 1353 2352 1358
rect 2708 1297 2714 1302
rect 2056 1253 2061 1258
rect 2100 1253 2105 1258
rect 2128 1255 2133 1260
rect 2127 1245 2132 1250
rect 2157 1253 2162 1258
rect 2535 1268 2541 1273
rect 2252 1149 2257 1154
rect 2282 1157 2287 1162
rect 2281 1147 2286 1152
rect 2309 1149 2314 1154
rect 2353 1149 2358 1154
rect 2551 1256 2556 1261
rect 2583 1256 2588 1261
rect 2708 1262 2714 1267
rect 2635 1256 2643 1261
rect 2496 1188 2501 1193
rect 2531 1187 2537 1192
rect 2470 1143 2475 1150
rect 2551 1140 2556 1145
rect 2613 1187 2619 1192
rect 2648 1186 2654 1191
rect 2584 1140 2589 1145
rect 2569 1129 2574 1135
rect 2673 1140 2681 1146
rect 2673 1094 2681 1103
rect 2255 1020 2260 1025
rect 2285 1028 2290 1033
rect 2284 1018 2289 1023
rect 2312 1020 2317 1025
rect 2356 1020 2361 1025
rect 2688 1003 2694 1008
rect 2858 1231 2864 1236
rect 2874 1219 2879 1224
rect 2906 1219 2911 1224
rect 2958 1219 2966 1224
rect 3097 1263 3103 1268
rect 2819 1151 2824 1156
rect 2854 1150 2860 1155
rect 2874 1103 2879 1108
rect 3113 1251 3118 1256
rect 3145 1251 3150 1256
rect 3197 1251 3205 1256
rect 3283 1251 3289 1262
rect 3058 1183 3063 1188
rect 3093 1182 3099 1187
rect 2936 1150 2942 1155
rect 2971 1149 2977 1154
rect 2907 1103 2912 1108
rect 2891 1093 2897 1099
rect 2996 1103 3004 1109
rect 3113 1135 3118 1140
rect 3175 1182 3181 1187
rect 3210 1181 3216 1186
rect 3146 1135 3151 1140
rect 3130 1126 3136 1131
rect 3235 1135 3243 1141
rect 3283 1168 3288 1173
rect 3355 1161 3360 1166
rect 3385 1169 3390 1174
rect 3384 1159 3389 1164
rect 3412 1161 3417 1166
rect 3456 1161 3461 1166
rect 2794 1043 2804 1049
rect 2865 1002 2870 1007
rect 2515 974 2521 979
rect 2531 962 2536 967
rect 2563 962 2568 967
rect 2688 968 2694 973
rect 2615 962 2623 967
rect 2476 894 2481 899
rect 2511 893 2517 898
rect 2265 859 2270 864
rect 2295 867 2300 872
rect 2294 857 2299 862
rect 2322 859 2327 864
rect 2366 859 2371 864
rect 2531 846 2536 851
rect 2593 893 2599 898
rect 2787 923 2792 929
rect 2628 892 2634 897
rect 2564 846 2569 851
rect 2549 835 2554 841
rect 2653 846 2661 852
rect 3291 1064 3296 1069
rect 3358 1025 3363 1030
rect 3388 1033 3393 1038
rect 3387 1023 3392 1028
rect 3415 1025 3420 1030
rect 3459 1025 3464 1030
rect 3383 860 3390 868
rect 2653 800 2661 809
rect 2838 792 2845 797
rect 2786 779 2791 784
rect 2853 779 2858 784
rect 2265 734 2270 739
rect 2295 742 2300 747
rect 2698 758 2704 763
rect 2294 732 2299 737
rect 2322 734 2327 739
rect 2366 734 2371 739
rect 2525 729 2531 734
rect 2541 717 2546 722
rect 2573 717 2578 722
rect 2698 723 2704 728
rect 2625 717 2633 722
rect 2486 649 2491 654
rect 2521 648 2527 653
rect 2541 601 2546 606
rect 2603 648 2609 653
rect 2865 700 2870 706
rect 3023 713 3029 719
rect 3082 702 3088 707
rect 2638 647 2644 652
rect 2574 601 2579 606
rect 2559 590 2564 596
rect 2663 601 2671 607
rect 3252 701 3258 708
rect 3236 681 3242 687
rect 3217 648 3227 653
rect 3236 602 3242 607
rect 2265 568 2270 573
rect 2295 576 2300 581
rect 3197 581 3206 589
rect 3383 578 3390 586
rect 2294 566 2299 571
rect 2322 568 2327 573
rect 2366 568 2371 573
rect 2853 570 2858 575
rect 2663 555 2671 564
rect 2797 558 2803 564
rect 2865 532 2870 537
rect 2713 504 2719 509
rect 2265 443 2270 448
rect 2295 451 2300 456
rect 2294 441 2299 446
rect 2322 443 2327 448
rect 2366 443 2371 448
rect 2540 475 2546 480
rect 2556 463 2561 468
rect 2588 463 2593 468
rect 2713 469 2719 474
rect 2640 463 2648 468
rect 3023 478 3029 484
rect 3176 480 3183 485
rect 3236 480 3242 486
rect 2501 395 2506 400
rect 2536 394 2542 399
rect 2556 347 2561 352
rect 2618 394 2624 399
rect 2838 453 2845 459
rect 3013 455 3019 460
rect 2653 393 2659 398
rect 2589 347 2594 352
rect 2574 336 2579 342
rect 2678 347 2686 353
rect 3218 415 3227 423
rect 2313 300 2318 305
rect 2343 308 2348 313
rect 2342 298 2347 303
rect 2370 300 2375 305
rect 2414 300 2419 305
rect 2678 301 2686 310
rect 3131 327 3136 333
rect 3144 327 3149 333
rect 3180 303 3188 309
rect 3280 290 3286 295
rect 3296 278 3301 283
rect 3328 278 3333 283
rect 3380 278 3388 283
rect 3241 210 3246 215
rect 3276 209 3282 214
rect 3296 162 3301 167
rect 3358 209 3364 214
rect 3393 208 3399 213
rect 3450 205 3456 211
rect 3329 162 3334 167
rect 3313 151 3319 158
rect 3418 162 3426 168
rect 3469 140 3474 145
rect 3501 132 3506 137
rect 3531 140 3536 145
rect 3530 130 3535 135
rect 3558 132 3563 137
rect 3602 132 3607 137
rect 2955 38 2960 43
rect 2985 46 2990 51
rect 2984 36 2989 41
rect 3012 38 3017 43
rect 3056 38 3061 43
<< metal2 >>
rect 2276 1411 2307 1414
rect 2276 1366 2280 1411
rect 2303 1358 2307 1411
rect 2225 1353 2246 1357
rect 2237 1329 2243 1353
rect 2276 1329 2280 1351
rect 2347 1329 2352 1353
rect 2237 1325 2356 1329
rect 2455 1315 2751 1316
rect 2455 1311 3289 1315
rect 2052 1282 2171 1286
rect 2056 1258 2061 1282
rect 2128 1260 2132 1282
rect 2165 1258 2171 1282
rect 2162 1254 2183 1258
rect 2101 1200 2105 1253
rect 2128 1200 2132 1245
rect 2101 1197 2132 1200
rect 2282 1207 2313 1210
rect 2282 1162 2286 1207
rect 2309 1154 2313 1207
rect 2231 1149 2252 1153
rect 2243 1125 2249 1149
rect 2282 1125 2286 1147
rect 2353 1125 2358 1149
rect 2243 1121 2362 1125
rect 2285 1078 2316 1081
rect 2285 1033 2289 1078
rect 2312 1025 2316 1078
rect 2234 1020 2255 1024
rect 2246 996 2252 1020
rect 2285 996 2289 1018
rect 2356 996 2361 1020
rect 2246 992 2365 996
rect 2295 917 2326 920
rect 2295 872 2299 917
rect 2322 864 2326 917
rect 2244 859 2265 863
rect 2256 835 2262 859
rect 2295 835 2299 857
rect 2366 835 2371 859
rect 2256 831 2375 835
rect 2295 792 2326 795
rect 2295 747 2299 792
rect 2322 739 2326 792
rect 2244 734 2265 738
rect 2256 710 2262 734
rect 2295 710 2299 732
rect 2366 710 2371 734
rect 2256 706 2375 710
rect 2295 626 2326 629
rect 2295 581 2299 626
rect 2322 573 2326 626
rect 2244 568 2265 572
rect 2256 544 2262 568
rect 2295 544 2299 566
rect 2366 544 2371 568
rect 2456 551 2461 1311
rect 2541 1268 2654 1273
rect 2496 1256 2551 1261
rect 2556 1256 2583 1261
rect 2588 1256 2635 1261
rect 2496 1193 2500 1256
rect 2531 1145 2537 1187
rect 2613 1146 2619 1187
rect 2648 1191 2654 1268
rect 2708 1267 2714 1297
rect 3103 1263 3216 1268
rect 3058 1251 3113 1256
rect 3118 1251 3145 1256
rect 3150 1251 3197 1256
rect 2864 1231 2977 1236
rect 2819 1219 2874 1224
rect 2879 1219 2906 1224
rect 2911 1219 2958 1224
rect 2819 1156 2823 1219
rect 2470 1114 2475 1143
rect 2530 1140 2551 1145
rect 2556 1140 2584 1145
rect 2589 1140 2603 1145
rect 2613 1140 2673 1146
rect 2569 1114 2574 1129
rect 2470 1107 2574 1114
rect 2673 1103 2681 1140
rect 2854 1108 2860 1150
rect 2936 1109 2942 1150
rect 2971 1154 2977 1231
rect 3058 1188 3062 1251
rect 3093 1140 3099 1182
rect 3175 1141 3181 1182
rect 3210 1186 3216 1263
rect 3283 1262 3289 1311
rect 3385 1219 3416 1222
rect 3385 1174 3389 1219
rect 3092 1135 3113 1140
rect 3118 1135 3146 1140
rect 3151 1135 3165 1140
rect 3175 1135 3235 1141
rect 2853 1103 2874 1108
rect 2879 1103 2907 1108
rect 2912 1103 2926 1108
rect 2936 1103 2996 1109
rect 3130 1107 3136 1126
rect 3283 1107 3288 1168
rect 3412 1166 3416 1219
rect 3334 1161 3355 1165
rect 3346 1137 3352 1161
rect 3385 1137 3389 1159
rect 3456 1137 3461 1161
rect 3346 1133 3465 1137
rect 3130 1102 3288 1107
rect 2891 1069 2897 1093
rect 3388 1083 3419 1086
rect 2891 1064 3291 1069
rect 2787 1043 2794 1049
rect 2521 974 2634 979
rect 2476 962 2531 967
rect 2536 962 2563 967
rect 2568 962 2615 967
rect 2476 899 2480 962
rect 2511 851 2517 893
rect 2593 852 2599 893
rect 2628 897 2634 974
rect 2688 973 2694 1003
rect 2787 929 2791 1043
rect 3388 1038 3392 1083
rect 3415 1030 3419 1083
rect 3337 1025 3358 1029
rect 2510 846 2531 851
rect 2536 846 2564 851
rect 2569 846 2583 851
rect 2593 846 2653 852
rect 2549 796 2554 835
rect 2653 809 2661 846
rect 2787 796 2791 923
rect 2549 789 2791 796
rect 2549 788 2554 789
rect 2531 729 2644 734
rect 2486 717 2541 722
rect 2546 717 2573 722
rect 2578 717 2625 722
rect 2486 654 2490 717
rect 2521 606 2527 648
rect 2603 607 2609 648
rect 2638 652 2644 729
rect 2698 728 2704 758
rect 2520 601 2541 606
rect 2546 601 2574 606
rect 2579 601 2593 606
rect 2603 601 2663 607
rect 2559 551 2564 590
rect 2663 564 2671 601
rect 2786 551 2790 779
rect 2456 545 2790 551
rect 2559 544 2790 545
rect 2256 540 2375 544
rect 2559 543 2564 544
rect 2295 501 2326 504
rect 2295 456 2299 501
rect 2322 448 2326 501
rect 2546 475 2659 480
rect 2501 463 2556 468
rect 2561 463 2588 468
rect 2593 463 2640 468
rect 2244 443 2265 447
rect 2256 419 2262 443
rect 2295 419 2299 441
rect 2366 419 2371 443
rect 2256 415 2375 419
rect 2501 400 2505 463
rect 2343 358 2374 361
rect 2343 313 2347 358
rect 2370 305 2374 358
rect 2536 352 2542 394
rect 2618 353 2624 394
rect 2653 398 2659 475
rect 2713 474 2719 504
rect 2535 347 2556 352
rect 2561 347 2589 352
rect 2594 347 2608 352
rect 2618 347 2678 353
rect 2292 300 2313 304
rect 2304 276 2310 300
rect 2343 276 2347 298
rect 2414 276 2419 300
rect 2574 297 2579 336
rect 2678 310 2686 347
rect 2797 297 2802 558
rect 2838 459 2845 792
rect 2853 575 2858 779
rect 2865 706 2870 1002
rect 3349 1001 3355 1025
rect 3388 1001 3392 1023
rect 3459 1001 3464 1025
rect 3349 997 3468 1001
rect 2865 537 2870 700
rect 3023 484 3029 713
rect 3082 661 3088 702
rect 3176 695 3258 701
rect 3176 661 3183 695
rect 3082 656 3183 661
rect 3218 653 3227 654
rect 3013 333 3019 455
rect 3176 355 3183 480
rect 3144 350 3183 355
rect 3144 333 3149 350
rect 3013 327 3131 333
rect 3197 309 3206 581
rect 3218 423 3227 648
rect 3236 607 3242 681
rect 3236 486 3242 602
rect 3383 586 3390 860
rect 3188 303 3206 309
rect 2574 290 2802 297
rect 3286 290 3399 295
rect 2574 289 2579 290
rect 2304 272 2423 276
rect 2797 129 2802 290
rect 3241 278 3296 283
rect 3301 278 3328 283
rect 3333 278 3380 283
rect 3241 215 3245 278
rect 3276 167 3282 209
rect 3358 168 3364 209
rect 3393 213 3399 290
rect 3456 205 3669 211
rect 3531 190 3562 193
rect 3275 162 3296 167
rect 3301 162 3329 167
rect 3334 162 3348 167
rect 3358 162 3418 168
rect 3319 151 3474 156
rect 3469 145 3474 151
rect 3531 145 3535 190
rect 3558 137 3562 190
rect 3480 132 3501 136
rect 2797 121 3450 129
rect 2797 113 2802 121
rect 2985 96 3016 99
rect 2985 51 2989 96
rect 3012 43 3016 96
rect 3444 86 3450 121
rect 3492 108 3498 132
rect 3531 108 3535 130
rect 3602 108 3607 132
rect 3492 104 3611 108
rect 3664 86 3669 205
rect 3444 81 3669 86
rect 2934 38 2955 42
rect 2946 14 2952 38
rect 2985 14 2989 36
rect 3056 14 3061 38
rect 2946 10 3065 14
<< m3contact >>
rect 2982 891 2988 897
rect 3215 860 3225 868
rect 2982 839 2988 845
rect 3215 811 3225 819
rect 2994 803 2999 809
rect 2994 768 2999 773
rect 2981 581 2988 589
rect 2981 518 2988 526
rect 3133 581 3139 589
rect 2867 328 2873 333
rect 2929 328 2935 333
<< m123contact >>
rect 3098 1026 3104 1031
rect 2982 1006 2987 1012
rect 2874 923 2879 929
rect 2982 925 2987 930
rect 3036 858 3043 864
rect 3076 839 3083 845
rect 3098 814 3104 819
rect 2874 792 2879 797
rect 3076 713 3083 719
rect 3036 648 3043 653
<< metal3 >>
rect 2982 930 2987 1006
rect 2874 797 2879 923
rect 2982 845 2988 891
rect 2994 773 2999 803
rect 3036 653 3043 858
rect 3076 719 3083 839
rect 3098 819 3104 1026
rect 3215 819 3225 860
rect 2981 526 2988 581
rect 3133 543 3139 581
rect 2873 328 2929 333
<< labels >>
rlabel metal1 2905 860 2958 864 1 Gnd
rlabel metal1 2905 860 2958 864 1 GND
rlabel metal1 2886 925 2905 927 1 P1
rlabel metal1 3011 893 3021 895 1 G1
rlabel metal1 3026 1028 3079 1032 5 VDD
rlabel metal1 2892 805 2945 809 5 VDD
rlabel metal1 2887 616 2940 620 1 Gnd
rlabel metal1 2887 616 2940 620 1 GND
rlabel metal1 3108 813 3161 817 5 VDD
rlabel metal1 2896 781 2912 783 1 P2
rlabel metal1 3141 893 3169 896 1 C2
rlabel metal1 3272 862 3325 866 5 VDD
rlabel metal1 3250 683 3268 685 1 G2
rlabel metal1 3350 683 3374 686 1 C3
rlabel metal1 2876 347 2929 351 1 Gnd
rlabel metal1 2876 347 2929 351 1 GND
rlabel metal1 2881 583 2934 587 5 VDD
rlabel metal1 3068 583 3121 587 5 VDD
rlabel metal1 3063 372 3116 376 1 Gnd
rlabel metal1 3063 372 3116 376 1 GND
rlabel metal1 2904 561 2925 563 1 P3
rlabel metal1 3292 580 3345 584 5 VDD
rlabel metal1 3287 417 3340 421 1 Gnd
rlabel metal1 3287 417 3340 421 1 GND
rlabel metal1 3182 236 3186 289 7 VDD
rlabel metal1 2885 241 2889 294 3 Gnd
rlabel metal1 2885 241 2889 294 3 GND
rlabel metal1 2931 303 2933 318 1 G3
rlabel metal1 3082 893 3089 895 1 C2
rlabel metal1 2571 987 2685 992 5 VDD
rlabel metal1 2595 827 2613 829 1 GND
rlabel metal1 2591 1281 2705 1286 5 VDD
rlabel metal1 2615 1121 2633 1123 1 GND
rlabel metal1 2581 742 2695 747 5 VDD
rlabel metal1 2605 582 2623 584 1 GND
rlabel metal1 2596 488 2710 493 5 VDD
rlabel metal1 2620 328 2638 330 1 GND
rlabel metal1 2751 892 2754 895 1 g1
rlabel metal1 2761 647 2764 650 1 g2
rlabel metal1 2776 393 2779 396 1 g3
rlabel metal1 2771 1186 2774 1189 1 C0
rlabel metal1 2910 1003 2929 1005 1 C0
rlabel metal1 2914 1244 3028 1249 5 VDD
rlabel metal1 2890 1082 3004 1088 1 GND
rlabel metal1 3153 1276 3267 1281 5 VDD
rlabel metal1 3129 1114 3243 1120 1 GND
rlabel metal1 3336 303 3450 308 5 VDD
rlabel metal1 3312 141 3426 147 1 GND
rlabel metal1 2255 1333 2258 1334 1 gnd
rlabel metal1 2261 1405 2263 1406 5 vdd
rlabel metal2 2240 1354 2244 1357 1 clk
rlabel metal1 2240 1362 2242 1364 1 a0
rlabel metal1 2261 1129 2264 1130 1 gnd
rlabel metal1 2267 1201 2269 1202 5 vdd
rlabel metal2 2246 1150 2250 1153 1 clk
rlabel metal1 2264 1000 2267 1001 1 gnd
rlabel metal1 2270 1072 2272 1073 5 vdd
rlabel metal2 2249 1021 2253 1024 1 clk
rlabel metal1 2274 839 2277 840 1 gnd
rlabel metal1 2280 911 2282 912 5 vdd
rlabel metal2 2259 860 2263 863 1 clk
rlabel metal1 2274 714 2277 715 1 gnd
rlabel metal1 2280 786 2282 787 5 vdd
rlabel metal2 2259 735 2263 738 1 clk
rlabel metal1 2274 548 2277 549 1 gnd
rlabel metal1 2280 620 2282 621 5 vdd
rlabel metal2 2259 569 2263 572 1 clk
rlabel metal1 2274 423 2277 424 1 gnd
rlabel metal1 2280 495 2282 496 5 vdd
rlabel metal2 2259 444 2263 447 1 clk
rlabel metal1 2246 1158 2248 1160 1 b0
rlabel metal1 2249 1029 2251 1031 1 a1
rlabel metal1 2259 868 2261 870 1 b1
rlabel metal1 2259 743 2261 745 1 a2
rlabel metal1 2259 577 2261 579 1 b2
rlabel metal1 2259 452 2261 454 1 a3
rlabel metal1 2322 280 2325 281 1 gnd
rlabel metal1 2328 352 2330 353 5 vdd
rlabel metal2 2307 301 2311 304 1 clk
rlabel metal1 2307 309 2309 311 1 b3
rlabel metal1 2150 1277 2153 1278 5 gnd
rlabel metal1 2145 1205 2147 1206 1 vdd
rlabel metal2 2164 1254 2168 1257 5 clk
rlabel metal1 3364 1141 3367 1142 1 gnd
rlabel metal1 3370 1213 3372 1214 5 vdd
rlabel metal2 3349 1162 3353 1165 1 clk
rlabel metal1 3349 1170 3351 1172 1 a0
rlabel metal1 3367 1005 3370 1006 1 gnd
rlabel metal1 3373 1077 3375 1078 5 vdd
rlabel metal2 3352 1026 3356 1029 1 clk
rlabel metal1 3352 1034 3354 1036 1 a0
rlabel metal1 2964 18 2967 19 1 gnd
rlabel metal1 2970 90 2972 91 5 vdd
rlabel metal2 2949 39 2953 42 1 clk
rlabel metal1 3510 112 3513 113 1 gnd
rlabel metal1 3516 184 3518 185 5 vdd
rlabel metal2 3495 133 3499 136 1 clk
rlabel metal1 2006 1295 2008 1297 3 sum0
rlabel metal1 3512 990 3514 993 1 sum1
rlabel metal1 3508 1124 3511 1128 1 sum2
rlabel metal1 3655 98 3657 100 7 sum3
rlabel metal1 3109 0 3111 3 1 C4
<< end >>
