magic
tech scmos
timestamp 1732097524
<< nwell >>
rect 1123 1041 1148 1098
rect 1160 1013 1185 1053
rect 1193 1046 1218 1086
rect 1236 1040 1261 1097
rect 1307 1039 1378 1102
rect 1446 1004 1471 1061
rect 1483 976 1508 1016
rect 1516 1009 1541 1049
rect 1559 1003 1584 1060
rect 1685 1036 1710 1093
rect 1722 1008 1747 1048
rect 1755 1041 1780 1081
rect 1798 1035 1823 1092
rect 1103 747 1128 804
rect 1140 719 1165 759
rect 1173 752 1198 792
rect 1216 746 1241 803
rect 1287 745 1358 808
rect 1522 779 1594 842
rect 1638 746 1710 847
rect 1113 502 1138 559
rect 1150 474 1175 514
rect 1183 507 1208 547
rect 1226 501 1251 558
rect 1297 500 1368 563
rect 1504 556 1571 619
rect 1589 611 1618 619
rect 1588 556 1618 611
rect 1720 569 1792 632
rect 1884 536 1976 681
rect 1493 309 1607 372
rect 1680 334 1747 397
rect 1765 334 1794 397
rect 1904 336 1976 399
rect 1128 248 1153 305
rect 1165 220 1190 260
rect 1198 253 1223 293
rect 1241 247 1266 304
rect 1312 246 1383 309
rect 1558 28 1744 142
rect 1868 63 1893 120
rect 1905 35 1930 75
rect 1938 68 1963 108
rect 1981 62 2006 119
rect 1558 25 1736 28
<< ntransistor >>
rect 1171 1063 1173 1083
rect 1134 1011 1136 1031
rect 1204 1016 1206 1036
rect 1247 1010 1249 1030
rect 1318 982 1320 1022
rect 1339 982 1341 1022
rect 1364 1009 1366 1029
rect 1494 1026 1496 1046
rect 1733 1058 1735 1078
rect 1457 974 1459 994
rect 1527 979 1529 999
rect 1696 1006 1698 1026
rect 1766 1011 1768 1031
rect 1809 1005 1811 1025
rect 1570 973 1572 993
rect 1151 769 1153 789
rect 1114 717 1116 737
rect 1184 722 1186 742
rect 1227 716 1229 736
rect 1298 688 1300 728
rect 1319 688 1321 728
rect 1344 715 1346 735
rect 1534 722 1536 762
rect 1555 722 1557 762
rect 1580 749 1582 769
rect 1650 714 1652 734
rect 1671 714 1673 734
rect 1696 716 1698 736
rect 1161 524 1163 544
rect 1124 472 1126 492
rect 1194 477 1196 497
rect 1237 471 1239 491
rect 1308 443 1310 483
rect 1329 443 1331 483
rect 1354 470 1356 490
rect 1516 479 1518 539
rect 1537 479 1539 539
rect 1558 479 1560 539
rect 1604 526 1606 546
rect 1732 512 1734 552
rect 1753 512 1755 552
rect 1778 539 1780 559
rect 1896 504 1898 524
rect 1917 504 1919 524
rect 1938 504 1940 524
rect 1962 506 1964 526
rect 1176 270 1178 290
rect 1139 218 1141 238
rect 1209 223 1211 243
rect 1252 217 1254 237
rect 1323 189 1325 229
rect 1344 189 1346 229
rect 1369 216 1371 236
rect 1505 212 1507 292
rect 1526 212 1528 292
rect 1547 212 1549 292
rect 1568 212 1570 292
rect 1593 279 1595 299
rect 1692 257 1694 317
rect 1713 257 1715 317
rect 1734 257 1736 317
rect 1780 304 1782 324
rect 1916 279 1918 319
rect 1937 279 1939 319
rect 1962 306 1964 326
rect 1521 128 1541 130
rect 1521 107 1541 109
rect 1521 86 1541 88
rect 1916 85 1918 105
rect 1521 65 1541 67
rect 1528 40 1548 42
rect 1879 33 1881 53
rect 1949 38 1951 58
rect 1992 32 1994 52
<< ptransistor >>
rect 1134 1051 1136 1091
rect 1204 1056 1206 1076
rect 1247 1050 1249 1090
rect 1171 1023 1173 1043
rect 1318 1049 1320 1089
rect 1339 1049 1341 1089
rect 1364 1049 1366 1089
rect 1457 1014 1459 1054
rect 1527 1019 1529 1039
rect 1570 1013 1572 1053
rect 1696 1046 1698 1086
rect 1766 1051 1768 1071
rect 1809 1045 1811 1085
rect 1494 986 1496 1006
rect 1733 1018 1735 1038
rect 1114 757 1116 797
rect 1184 762 1186 782
rect 1227 756 1229 796
rect 1151 729 1153 749
rect 1298 755 1300 795
rect 1319 755 1321 795
rect 1344 755 1346 795
rect 1534 789 1536 829
rect 1555 789 1557 829
rect 1580 789 1582 829
rect 1650 756 1652 836
rect 1671 756 1673 836
rect 1696 756 1698 796
rect 1124 512 1126 552
rect 1194 517 1196 537
rect 1237 511 1239 551
rect 1516 566 1518 606
rect 1537 566 1539 606
rect 1558 566 1560 606
rect 1604 566 1606 606
rect 1732 579 1734 619
rect 1753 579 1755 619
rect 1778 579 1780 619
rect 1161 484 1163 504
rect 1308 510 1310 550
rect 1329 510 1331 550
rect 1354 510 1356 550
rect 1896 545 1898 665
rect 1917 545 1919 665
rect 1938 545 1940 665
rect 1962 546 1964 586
rect 1505 319 1507 359
rect 1526 319 1528 359
rect 1547 319 1549 359
rect 1568 319 1570 359
rect 1593 319 1595 359
rect 1692 344 1694 384
rect 1713 344 1715 384
rect 1734 344 1736 384
rect 1780 344 1782 384
rect 1916 346 1918 386
rect 1937 346 1939 386
rect 1962 346 1964 386
rect 1139 258 1141 298
rect 1209 263 1211 283
rect 1252 257 1254 297
rect 1176 230 1178 250
rect 1323 256 1325 296
rect 1344 256 1346 296
rect 1369 256 1371 296
rect 1568 128 1728 130
rect 1568 107 1728 109
rect 1568 86 1728 88
rect 1879 73 1881 113
rect 1949 78 1951 98
rect 1568 65 1728 67
rect 1992 72 1994 112
rect 1568 40 1608 42
rect 1916 45 1918 65
<< ndiffusion >>
rect 1170 1063 1171 1083
rect 1173 1063 1174 1083
rect 1133 1011 1134 1031
rect 1136 1011 1137 1031
rect 1203 1016 1204 1036
rect 1206 1016 1207 1036
rect 1246 1010 1247 1030
rect 1249 1010 1250 1030
rect 1317 982 1318 1022
rect 1320 982 1321 1022
rect 1338 982 1339 1022
rect 1341 982 1342 1022
rect 1363 1009 1364 1029
rect 1366 1009 1367 1029
rect 1493 1026 1494 1046
rect 1496 1026 1497 1046
rect 1732 1058 1733 1078
rect 1735 1058 1736 1078
rect 1456 974 1457 994
rect 1459 974 1460 994
rect 1526 979 1527 999
rect 1529 979 1530 999
rect 1695 1006 1696 1026
rect 1698 1006 1699 1026
rect 1765 1011 1766 1031
rect 1768 1011 1769 1031
rect 1808 1005 1809 1025
rect 1811 1005 1812 1025
rect 1569 973 1570 993
rect 1572 973 1573 993
rect 1150 769 1151 789
rect 1153 769 1154 789
rect 1113 717 1114 737
rect 1116 717 1117 737
rect 1183 722 1184 742
rect 1186 722 1187 742
rect 1226 716 1227 736
rect 1229 716 1230 736
rect 1297 688 1298 728
rect 1300 688 1301 728
rect 1318 688 1319 728
rect 1321 688 1322 728
rect 1343 715 1344 735
rect 1346 715 1347 735
rect 1533 722 1534 762
rect 1536 722 1537 762
rect 1554 722 1555 762
rect 1557 722 1558 762
rect 1579 749 1580 769
rect 1582 749 1583 769
rect 1649 714 1650 734
rect 1652 714 1653 734
rect 1670 714 1671 734
rect 1673 714 1674 734
rect 1695 716 1696 736
rect 1698 716 1699 736
rect 1160 524 1161 544
rect 1163 524 1164 544
rect 1123 472 1124 492
rect 1126 472 1127 492
rect 1193 477 1194 497
rect 1196 477 1197 497
rect 1236 471 1237 491
rect 1239 471 1240 491
rect 1307 443 1308 483
rect 1310 443 1311 483
rect 1328 443 1329 483
rect 1331 443 1332 483
rect 1353 470 1354 490
rect 1356 470 1357 490
rect 1515 479 1516 539
rect 1518 479 1519 539
rect 1536 479 1537 539
rect 1539 479 1540 539
rect 1557 479 1558 539
rect 1560 479 1561 539
rect 1603 526 1604 546
rect 1606 526 1607 546
rect 1731 512 1732 552
rect 1734 512 1735 552
rect 1752 512 1753 552
rect 1755 512 1756 552
rect 1777 539 1778 559
rect 1780 539 1781 559
rect 1895 504 1896 524
rect 1898 504 1899 524
rect 1916 504 1917 524
rect 1919 504 1920 524
rect 1937 504 1938 524
rect 1940 504 1941 524
rect 1961 506 1962 526
rect 1964 506 1965 526
rect 1175 270 1176 290
rect 1178 270 1179 290
rect 1138 218 1139 238
rect 1141 218 1142 238
rect 1208 223 1209 243
rect 1211 223 1212 243
rect 1251 217 1252 237
rect 1254 217 1255 237
rect 1322 189 1323 229
rect 1325 189 1326 229
rect 1343 189 1344 229
rect 1346 189 1347 229
rect 1368 216 1369 236
rect 1371 216 1372 236
rect 1504 212 1505 292
rect 1507 212 1508 292
rect 1525 212 1526 292
rect 1528 212 1529 292
rect 1546 212 1547 292
rect 1549 212 1550 292
rect 1567 212 1568 292
rect 1570 212 1571 292
rect 1592 279 1593 299
rect 1595 279 1596 299
rect 1691 257 1692 317
rect 1694 257 1695 317
rect 1712 257 1713 317
rect 1715 257 1716 317
rect 1733 257 1734 317
rect 1736 257 1737 317
rect 1779 304 1780 324
rect 1782 304 1783 324
rect 1915 279 1916 319
rect 1918 279 1919 319
rect 1936 279 1937 319
rect 1939 279 1940 319
rect 1961 306 1962 326
rect 1964 306 1965 326
rect 1521 130 1541 131
rect 1521 127 1541 128
rect 1521 109 1541 110
rect 1521 106 1541 107
rect 1521 88 1541 89
rect 1521 85 1541 86
rect 1915 85 1916 105
rect 1918 85 1919 105
rect 1521 67 1541 68
rect 1521 64 1541 65
rect 1528 42 1548 43
rect 1528 39 1548 40
rect 1878 33 1879 53
rect 1881 33 1882 53
rect 1948 38 1949 58
rect 1951 38 1952 58
rect 1991 32 1992 52
rect 1994 32 1995 52
<< pdiffusion >>
rect 1133 1051 1134 1091
rect 1136 1051 1137 1091
rect 1203 1056 1204 1076
rect 1206 1056 1207 1076
rect 1246 1050 1247 1090
rect 1249 1050 1250 1090
rect 1170 1023 1171 1043
rect 1173 1023 1174 1043
rect 1317 1049 1318 1089
rect 1320 1049 1321 1089
rect 1338 1049 1339 1089
rect 1341 1049 1342 1089
rect 1363 1049 1364 1089
rect 1366 1049 1367 1089
rect 1456 1014 1457 1054
rect 1459 1014 1460 1054
rect 1526 1019 1527 1039
rect 1529 1019 1530 1039
rect 1569 1013 1570 1053
rect 1572 1013 1573 1053
rect 1695 1046 1696 1086
rect 1698 1046 1699 1086
rect 1765 1051 1766 1071
rect 1768 1051 1769 1071
rect 1808 1045 1809 1085
rect 1811 1045 1812 1085
rect 1493 986 1494 1006
rect 1496 986 1497 1006
rect 1732 1018 1733 1038
rect 1735 1018 1736 1038
rect 1113 757 1114 797
rect 1116 757 1117 797
rect 1183 762 1184 782
rect 1186 762 1187 782
rect 1226 756 1227 796
rect 1229 756 1230 796
rect 1150 729 1151 749
rect 1153 729 1154 749
rect 1297 755 1298 795
rect 1300 755 1301 795
rect 1318 755 1319 795
rect 1321 755 1322 795
rect 1343 755 1344 795
rect 1346 755 1347 795
rect 1533 789 1534 829
rect 1536 789 1537 829
rect 1554 789 1555 829
rect 1557 789 1558 829
rect 1579 789 1580 829
rect 1582 789 1583 829
rect 1649 756 1650 836
rect 1652 756 1653 836
rect 1670 756 1671 836
rect 1673 756 1674 836
rect 1695 756 1696 796
rect 1698 756 1699 796
rect 1123 512 1124 552
rect 1126 512 1127 552
rect 1193 517 1194 537
rect 1196 517 1197 537
rect 1236 511 1237 551
rect 1239 511 1240 551
rect 1515 566 1516 606
rect 1518 566 1519 606
rect 1536 566 1537 606
rect 1539 566 1540 606
rect 1557 566 1558 606
rect 1560 566 1561 606
rect 1603 566 1604 606
rect 1606 566 1607 606
rect 1731 579 1732 619
rect 1734 579 1735 619
rect 1752 579 1753 619
rect 1755 579 1756 619
rect 1777 579 1778 619
rect 1780 579 1781 619
rect 1160 484 1161 504
rect 1163 484 1164 504
rect 1307 510 1308 550
rect 1310 510 1311 550
rect 1328 510 1329 550
rect 1331 510 1332 550
rect 1353 510 1354 550
rect 1356 510 1357 550
rect 1895 545 1896 665
rect 1898 545 1899 665
rect 1916 545 1917 665
rect 1919 545 1920 665
rect 1937 545 1938 665
rect 1940 545 1941 665
rect 1961 546 1962 586
rect 1964 546 1965 586
rect 1504 319 1505 359
rect 1507 319 1508 359
rect 1525 319 1526 359
rect 1528 319 1529 359
rect 1546 319 1547 359
rect 1549 319 1550 359
rect 1567 319 1568 359
rect 1570 319 1571 359
rect 1592 319 1593 359
rect 1595 319 1596 359
rect 1691 344 1692 384
rect 1694 344 1695 384
rect 1712 344 1713 384
rect 1715 344 1716 384
rect 1733 344 1734 384
rect 1736 344 1737 384
rect 1779 344 1780 384
rect 1782 344 1783 384
rect 1915 346 1916 386
rect 1918 346 1919 386
rect 1936 346 1937 386
rect 1939 346 1940 386
rect 1961 346 1962 386
rect 1964 346 1965 386
rect 1138 258 1139 298
rect 1141 258 1142 298
rect 1208 263 1209 283
rect 1211 263 1212 283
rect 1251 257 1252 297
rect 1254 257 1255 297
rect 1175 230 1176 250
rect 1178 230 1179 250
rect 1322 256 1323 296
rect 1325 256 1326 296
rect 1343 256 1344 296
rect 1346 256 1347 296
rect 1368 256 1369 296
rect 1371 256 1372 296
rect 1568 130 1728 131
rect 1568 127 1728 128
rect 1568 109 1728 110
rect 1568 106 1728 107
rect 1568 88 1728 89
rect 1568 85 1728 86
rect 1878 73 1879 113
rect 1881 73 1882 113
rect 1948 78 1949 98
rect 1951 78 1952 98
rect 1568 67 1728 68
rect 1568 64 1728 65
rect 1991 72 1992 112
rect 1994 72 1995 112
rect 1568 42 1608 43
rect 1568 39 1608 40
rect 1915 45 1916 65
rect 1918 45 1919 65
<< ndcontact >>
rect 1166 1063 1170 1083
rect 1174 1063 1178 1083
rect 1129 1011 1133 1031
rect 1137 1011 1141 1031
rect 1199 1016 1203 1036
rect 1207 1016 1211 1036
rect 1242 1010 1246 1030
rect 1250 1010 1254 1030
rect 1313 982 1317 1022
rect 1321 982 1338 1022
rect 1342 982 1346 1022
rect 1359 1009 1363 1029
rect 1367 1009 1371 1029
rect 1489 1026 1493 1046
rect 1497 1026 1501 1046
rect 1728 1058 1732 1078
rect 1736 1058 1740 1078
rect 1452 974 1456 994
rect 1460 974 1464 994
rect 1522 979 1526 999
rect 1530 979 1534 999
rect 1691 1006 1695 1026
rect 1699 1006 1703 1026
rect 1761 1011 1765 1031
rect 1769 1011 1773 1031
rect 1804 1005 1808 1025
rect 1812 1005 1816 1025
rect 1565 973 1569 993
rect 1573 973 1577 993
rect 1146 769 1150 789
rect 1154 769 1158 789
rect 1109 717 1113 737
rect 1117 717 1121 737
rect 1179 722 1183 742
rect 1187 722 1191 742
rect 1222 716 1226 736
rect 1230 716 1234 736
rect 1293 688 1297 728
rect 1301 688 1318 728
rect 1322 688 1326 728
rect 1339 715 1343 735
rect 1347 715 1351 735
rect 1529 722 1533 762
rect 1537 722 1554 762
rect 1558 722 1562 762
rect 1575 749 1579 769
rect 1583 749 1587 769
rect 1645 714 1649 734
rect 1653 714 1657 734
rect 1666 714 1670 734
rect 1674 714 1678 734
rect 1691 716 1695 736
rect 1699 716 1703 736
rect 1156 524 1160 544
rect 1164 524 1168 544
rect 1119 472 1123 492
rect 1127 472 1131 492
rect 1189 477 1193 497
rect 1197 477 1201 497
rect 1232 471 1236 491
rect 1240 471 1244 491
rect 1303 443 1307 483
rect 1311 443 1328 483
rect 1332 443 1336 483
rect 1349 470 1353 490
rect 1357 470 1361 490
rect 1511 479 1515 539
rect 1519 479 1523 539
rect 1532 479 1536 539
rect 1540 479 1544 539
rect 1553 479 1557 539
rect 1561 479 1565 539
rect 1599 526 1603 546
rect 1607 526 1611 546
rect 1727 512 1731 552
rect 1735 512 1752 552
rect 1756 512 1760 552
rect 1773 539 1777 559
rect 1781 539 1785 559
rect 1891 504 1895 524
rect 1899 504 1903 524
rect 1912 504 1916 524
rect 1920 504 1924 524
rect 1933 504 1937 524
rect 1941 504 1945 524
rect 1957 506 1961 526
rect 1965 506 1969 526
rect 1171 270 1175 290
rect 1179 270 1183 290
rect 1134 218 1138 238
rect 1142 218 1146 238
rect 1204 223 1208 243
rect 1212 223 1216 243
rect 1247 217 1251 237
rect 1255 217 1259 237
rect 1318 189 1322 229
rect 1326 189 1343 229
rect 1347 189 1351 229
rect 1364 216 1368 236
rect 1372 216 1376 236
rect 1500 212 1504 292
rect 1508 212 1512 292
rect 1521 212 1525 292
rect 1529 212 1533 292
rect 1542 212 1546 292
rect 1550 212 1554 292
rect 1563 212 1567 292
rect 1571 212 1575 292
rect 1588 279 1592 299
rect 1596 279 1600 299
rect 1687 257 1691 317
rect 1695 257 1699 317
rect 1708 257 1712 317
rect 1716 257 1720 317
rect 1729 257 1733 317
rect 1737 257 1741 317
rect 1775 304 1779 324
rect 1783 304 1787 324
rect 1911 279 1915 319
rect 1919 279 1936 319
rect 1940 279 1944 319
rect 1957 306 1961 326
rect 1965 306 1969 326
rect 1521 131 1541 135
rect 1521 123 1541 127
rect 1521 110 1541 114
rect 1521 102 1541 106
rect 1521 89 1541 93
rect 1521 81 1541 85
rect 1911 85 1915 105
rect 1919 85 1923 105
rect 1521 68 1541 72
rect 1521 60 1541 64
rect 1528 43 1548 47
rect 1528 35 1548 39
rect 1874 33 1878 53
rect 1882 33 1886 53
rect 1944 38 1948 58
rect 1952 38 1956 58
rect 1987 32 1991 52
rect 1995 32 1999 52
<< pdcontact >>
rect 1129 1051 1133 1091
rect 1137 1051 1141 1091
rect 1199 1056 1203 1076
rect 1207 1056 1211 1076
rect 1242 1050 1246 1090
rect 1250 1050 1254 1090
rect 1166 1023 1170 1043
rect 1174 1023 1178 1043
rect 1313 1049 1317 1089
rect 1321 1049 1338 1089
rect 1342 1049 1346 1089
rect 1359 1049 1363 1089
rect 1367 1049 1371 1089
rect 1452 1014 1456 1054
rect 1460 1014 1464 1054
rect 1522 1019 1526 1039
rect 1530 1019 1534 1039
rect 1565 1013 1569 1053
rect 1573 1013 1577 1053
rect 1691 1046 1695 1086
rect 1699 1046 1703 1086
rect 1761 1051 1765 1071
rect 1769 1051 1773 1071
rect 1804 1045 1808 1085
rect 1812 1045 1816 1085
rect 1489 986 1493 1006
rect 1497 986 1501 1006
rect 1728 1018 1732 1038
rect 1736 1018 1740 1038
rect 1109 757 1113 797
rect 1117 757 1121 797
rect 1179 762 1183 782
rect 1187 762 1191 782
rect 1222 756 1226 796
rect 1230 756 1234 796
rect 1146 729 1150 749
rect 1154 729 1158 749
rect 1293 755 1297 795
rect 1301 755 1318 795
rect 1322 755 1326 795
rect 1339 755 1343 795
rect 1347 755 1351 795
rect 1529 789 1533 829
rect 1537 789 1554 829
rect 1558 789 1562 829
rect 1575 789 1579 829
rect 1583 789 1587 829
rect 1645 756 1649 836
rect 1653 756 1657 836
rect 1666 756 1670 836
rect 1674 756 1678 836
rect 1691 756 1695 796
rect 1699 756 1703 796
rect 1119 512 1123 552
rect 1127 512 1131 552
rect 1189 517 1193 537
rect 1197 517 1201 537
rect 1232 511 1236 551
rect 1240 511 1244 551
rect 1511 566 1515 606
rect 1519 566 1536 606
rect 1540 566 1557 606
rect 1561 566 1565 606
rect 1599 566 1603 606
rect 1607 566 1611 606
rect 1727 579 1731 619
rect 1735 579 1752 619
rect 1756 579 1760 619
rect 1773 579 1777 619
rect 1781 579 1785 619
rect 1156 484 1160 504
rect 1164 484 1168 504
rect 1303 510 1307 550
rect 1311 510 1328 550
rect 1332 510 1336 550
rect 1349 510 1353 550
rect 1357 510 1361 550
rect 1891 545 1895 665
rect 1899 545 1903 665
rect 1912 545 1916 665
rect 1920 545 1924 665
rect 1933 545 1937 665
rect 1941 545 1945 665
rect 1957 546 1961 586
rect 1965 546 1969 586
rect 1500 319 1504 359
rect 1508 319 1525 359
rect 1529 319 1546 359
rect 1550 319 1567 359
rect 1571 319 1575 359
rect 1588 319 1592 359
rect 1596 319 1600 359
rect 1687 344 1691 384
rect 1695 344 1712 384
rect 1716 344 1733 384
rect 1737 344 1741 384
rect 1775 344 1779 384
rect 1783 344 1787 384
rect 1911 346 1915 386
rect 1919 346 1936 386
rect 1940 346 1944 386
rect 1957 346 1961 386
rect 1965 346 1969 386
rect 1134 258 1138 298
rect 1142 258 1146 298
rect 1204 263 1208 283
rect 1212 263 1216 283
rect 1247 257 1251 297
rect 1255 257 1259 297
rect 1171 230 1175 250
rect 1179 230 1183 250
rect 1318 256 1322 296
rect 1326 256 1343 296
rect 1347 256 1351 296
rect 1364 256 1368 296
rect 1372 256 1376 296
rect 1568 131 1728 135
rect 1568 123 1728 127
rect 1568 110 1728 114
rect 1568 102 1728 106
rect 1568 89 1728 93
rect 1568 81 1728 85
rect 1874 73 1878 113
rect 1882 73 1886 113
rect 1944 78 1948 98
rect 1952 78 1956 98
rect 1568 68 1728 72
rect 1568 60 1728 64
rect 1987 72 1991 112
rect 1995 72 1999 112
rect 1568 43 1608 47
rect 1568 35 1608 39
rect 1911 45 1915 65
rect 1919 45 1923 65
<< polysilicon >>
rect 1134 1091 1136 1095
rect 1247 1090 1249 1094
rect 1171 1083 1173 1090
rect 1204 1076 1206 1090
rect 1171 1060 1173 1063
rect 1204 1053 1206 1056
rect 1134 1031 1136 1051
rect 1318 1089 1320 1093
rect 1339 1089 1341 1108
rect 1364 1089 1366 1093
rect 1171 1043 1173 1046
rect 1204 1036 1206 1039
rect 1134 1008 1136 1011
rect 1171 1009 1173 1023
rect 1247 1030 1249 1050
rect 1696 1086 1698 1090
rect 1457 1054 1459 1058
rect 1204 1009 1206 1016
rect 1318 1022 1320 1049
rect 1339 1022 1341 1049
rect 1364 1029 1366 1049
rect 1247 1007 1249 1010
rect 1570 1053 1572 1057
rect 1494 1046 1496 1053
rect 1527 1039 1529 1053
rect 1494 1023 1496 1026
rect 1527 1016 1529 1019
rect 1364 1006 1366 1009
rect 1457 994 1459 1014
rect 1809 1085 1811 1089
rect 1733 1078 1735 1085
rect 1766 1071 1768 1085
rect 1733 1055 1735 1058
rect 1766 1048 1768 1051
rect 1696 1026 1698 1046
rect 1733 1038 1735 1041
rect 1494 1006 1496 1009
rect 1318 979 1320 982
rect 1339 979 1341 982
rect 1527 999 1529 1002
rect 1457 971 1459 974
rect 1494 972 1496 986
rect 1570 993 1572 1013
rect 1766 1031 1768 1034
rect 1696 1003 1698 1006
rect 1733 1004 1735 1018
rect 1809 1025 1811 1045
rect 1766 1004 1768 1011
rect 1809 1002 1811 1005
rect 1527 972 1529 979
rect 1570 970 1572 973
rect 1534 829 1536 833
rect 1555 829 1557 848
rect 1650 836 1652 839
rect 1671 836 1673 853
rect 1580 829 1582 833
rect 1114 797 1116 801
rect 1227 796 1229 800
rect 1151 789 1153 796
rect 1184 782 1186 796
rect 1151 766 1153 769
rect 1184 759 1186 762
rect 1114 737 1116 757
rect 1298 795 1300 799
rect 1319 795 1321 814
rect 1344 795 1346 799
rect 1151 749 1153 752
rect 1184 742 1186 745
rect 1114 714 1116 717
rect 1151 715 1153 729
rect 1227 736 1229 756
rect 1534 762 1536 789
rect 1555 762 1557 789
rect 1580 769 1582 789
rect 1184 715 1186 722
rect 1298 728 1300 755
rect 1319 728 1321 755
rect 1344 735 1346 755
rect 1227 713 1229 716
rect 1696 796 1698 800
rect 1580 746 1582 749
rect 1650 734 1652 756
rect 1671 734 1673 756
rect 1696 736 1698 756
rect 1534 719 1536 722
rect 1555 719 1557 722
rect 1344 712 1346 715
rect 1650 711 1652 714
rect 1671 711 1673 714
rect 1696 713 1698 716
rect 1298 685 1300 688
rect 1319 685 1321 688
rect 1896 665 1898 673
rect 1917 665 1919 687
rect 1938 665 1940 697
rect 1516 606 1518 610
rect 1537 606 1539 625
rect 1558 606 1560 638
rect 1732 619 1734 623
rect 1753 619 1755 638
rect 1778 619 1780 623
rect 1604 606 1606 610
rect 1124 552 1126 556
rect 1237 551 1239 555
rect 1161 544 1163 551
rect 1194 537 1196 551
rect 1161 521 1163 524
rect 1194 514 1196 517
rect 1124 492 1126 512
rect 1308 550 1310 554
rect 1329 550 1331 569
rect 1354 550 1356 554
rect 1161 504 1163 507
rect 1194 497 1196 500
rect 1124 469 1126 472
rect 1161 470 1163 484
rect 1237 491 1239 511
rect 1516 539 1518 566
rect 1537 539 1539 566
rect 1558 539 1560 566
rect 1604 546 1606 566
rect 1732 552 1734 579
rect 1753 552 1755 579
rect 1778 559 1780 579
rect 1194 470 1196 477
rect 1308 483 1310 510
rect 1329 483 1331 510
rect 1354 490 1356 510
rect 1237 468 1239 471
rect 1604 523 1606 526
rect 1962 586 1964 590
rect 1778 536 1780 539
rect 1896 524 1898 545
rect 1917 524 1919 545
rect 1938 524 1940 545
rect 1962 526 1964 546
rect 1732 509 1734 512
rect 1753 509 1755 512
rect 1896 501 1898 504
rect 1917 501 1919 504
rect 1938 501 1940 504
rect 1962 503 1964 506
rect 1516 475 1518 479
rect 1537 475 1539 479
rect 1558 475 1560 479
rect 1354 467 1356 470
rect 1308 440 1310 443
rect 1329 440 1331 443
rect 1505 359 1507 363
rect 1526 359 1528 378
rect 1547 359 1549 405
rect 1568 359 1570 416
rect 1692 384 1694 388
rect 1713 384 1715 405
rect 1734 384 1736 416
rect 1780 384 1782 388
rect 1916 386 1918 390
rect 1937 386 1939 405
rect 1962 386 1964 390
rect 1593 359 1595 363
rect 1139 298 1141 302
rect 1252 297 1254 301
rect 1176 290 1178 297
rect 1209 283 1211 297
rect 1176 267 1178 270
rect 1209 260 1211 263
rect 1139 238 1141 258
rect 1323 296 1325 300
rect 1344 296 1346 315
rect 1369 296 1371 300
rect 1176 250 1178 253
rect 1209 243 1211 246
rect 1139 215 1141 218
rect 1176 216 1178 230
rect 1252 237 1254 257
rect 1505 292 1507 319
rect 1526 292 1528 319
rect 1547 292 1549 319
rect 1568 292 1570 319
rect 1593 299 1595 319
rect 1692 317 1694 344
rect 1713 317 1715 344
rect 1734 317 1736 344
rect 1780 324 1782 344
rect 1209 216 1211 223
rect 1323 229 1325 256
rect 1344 229 1346 256
rect 1369 236 1371 256
rect 1252 214 1254 217
rect 1369 213 1371 216
rect 1593 276 1595 279
rect 1916 319 1918 346
rect 1937 319 1939 346
rect 1962 326 1964 346
rect 1780 301 1782 304
rect 1962 303 1964 306
rect 1916 276 1918 279
rect 1937 276 1939 279
rect 1692 253 1694 257
rect 1713 253 1715 257
rect 1734 253 1736 257
rect 1505 209 1507 212
rect 1526 209 1528 212
rect 1547 209 1549 212
rect 1568 209 1570 212
rect 1323 186 1325 189
rect 1344 186 1346 189
rect 1517 128 1521 130
rect 1541 128 1568 130
rect 1728 128 1735 130
rect 1879 113 1881 117
rect 1517 107 1521 109
rect 1541 107 1568 109
rect 1728 107 1750 109
rect 1517 86 1521 88
rect 1541 86 1568 88
rect 1728 86 1763 88
rect 1992 112 1994 116
rect 1916 105 1918 112
rect 1949 98 1951 112
rect 1916 82 1918 85
rect 1949 75 1951 78
rect 1517 65 1521 67
rect 1541 65 1568 67
rect 1728 65 1774 67
rect 1879 53 1881 73
rect 1916 65 1918 68
rect 1525 40 1528 42
rect 1548 40 1568 42
rect 1608 40 1735 42
rect 1949 58 1951 61
rect 1879 30 1881 33
rect 1916 31 1918 45
rect 1992 52 1994 72
rect 1949 31 1951 38
rect 1992 29 1994 32
<< polycontact >>
rect 1337 1108 1343 1113
rect 1170 1090 1174 1095
rect 1203 1090 1207 1095
rect 1130 1034 1134 1039
rect 1243 1033 1247 1038
rect 1311 1029 1318 1035
rect 1360 1032 1364 1037
rect 1170 1004 1174 1009
rect 1203 1004 1207 1009
rect 1493 1053 1497 1058
rect 1526 1053 1530 1058
rect 1453 997 1457 1002
rect 1732 1085 1736 1090
rect 1765 1085 1769 1090
rect 1692 1029 1696 1034
rect 1566 996 1570 1001
rect 1805 1028 1809 1033
rect 1732 999 1736 1004
rect 1765 999 1769 1004
rect 1493 967 1497 972
rect 1526 967 1530 972
rect 1669 853 1675 858
rect 1553 848 1559 853
rect 1317 814 1323 819
rect 1150 796 1154 801
rect 1183 796 1187 801
rect 1110 740 1114 745
rect 1223 739 1227 744
rect 1527 769 1534 775
rect 1576 772 1580 777
rect 1291 735 1298 741
rect 1340 738 1344 743
rect 1150 710 1154 715
rect 1183 710 1187 715
rect 1643 737 1650 743
rect 1692 739 1696 744
rect 1936 697 1942 702
rect 1915 687 1921 692
rect 1556 638 1562 643
rect 1751 638 1757 643
rect 1535 625 1541 630
rect 1327 569 1333 574
rect 1160 551 1164 556
rect 1193 551 1197 556
rect 1120 495 1124 500
rect 1233 494 1237 499
rect 1509 546 1516 552
rect 1600 549 1604 554
rect 1725 559 1732 565
rect 1774 562 1778 567
rect 1301 490 1308 496
rect 1350 493 1354 498
rect 1160 465 1164 470
rect 1193 465 1197 470
rect 1889 527 1896 533
rect 1958 529 1962 534
rect 1566 416 1572 421
rect 1732 416 1738 421
rect 1545 405 1551 410
rect 1524 378 1530 383
rect 1711 405 1717 410
rect 1935 405 1941 410
rect 1342 315 1348 320
rect 1685 324 1692 330
rect 1175 297 1179 302
rect 1208 297 1212 302
rect 1135 241 1139 246
rect 1498 299 1505 305
rect 1248 240 1252 245
rect 1589 302 1593 307
rect 1776 327 1780 332
rect 1909 326 1916 332
rect 1316 236 1323 242
rect 1365 239 1369 244
rect 1175 211 1179 216
rect 1208 211 1212 216
rect 1958 329 1962 334
rect 1548 130 1554 137
rect 1750 105 1755 111
rect 1763 84 1768 90
rect 1915 112 1919 117
rect 1948 112 1952 117
rect 1774 63 1779 69
rect 1875 56 1879 61
rect 1551 42 1556 46
rect 1988 55 1992 60
rect 1915 26 1919 31
rect 1948 26 1952 31
<< metal1 >>
rect 1321 1143 1327 1148
rect 1114 1127 1376 1132
rect 1129 1091 1133 1127
rect 1154 1059 1159 1114
rect 1170 1095 1174 1102
rect 1203 1095 1207 1102
rect 1242 1090 1246 1127
rect 1289 1108 1327 1113
rect 1333 1108 1337 1113
rect 1343 1108 1345 1113
rect 1289 1107 1300 1108
rect 1262 1102 1300 1107
rect 1370 1102 1376 1127
rect 1663 1122 1896 1127
rect 1307 1094 1378 1102
rect 1396 1100 1667 1105
rect 1166 1059 1170 1063
rect 1154 1055 1170 1059
rect 1120 1034 1130 1039
rect 1137 1038 1141 1051
rect 1166 1043 1170 1055
rect 1137 1033 1150 1038
rect 1137 1031 1141 1033
rect 1174 1058 1178 1063
rect 1174 1054 1192 1058
rect 1174 1043 1178 1054
rect 1187 1044 1192 1054
rect 1199 1044 1203 1056
rect 1187 1040 1203 1044
rect 1188 1039 1203 1040
rect 1129 972 1133 1011
rect 1170 991 1174 1004
rect 1188 981 1193 1039
rect 1199 1036 1203 1039
rect 1207 1043 1211 1056
rect 1207 1039 1228 1043
rect 1207 1036 1211 1039
rect 1222 1038 1228 1039
rect 1222 1033 1232 1038
rect 1238 1033 1243 1038
rect 1250 1037 1254 1050
rect 1313 1089 1317 1094
rect 1342 1089 1346 1094
rect 1359 1089 1363 1094
rect 1250 1032 1267 1037
rect 1250 1030 1254 1032
rect 1292 1029 1311 1035
rect 1326 1030 1331 1049
rect 1352 1032 1360 1037
rect 1367 1036 1371 1049
rect 1396 1036 1400 1100
rect 1424 1090 1657 1095
rect 1352 1030 1356 1032
rect 1203 991 1207 1004
rect 1242 972 1246 1010
rect 1292 992 1300 1029
rect 1326 1026 1356 1030
rect 1367 1031 1400 1036
rect 1367 1029 1371 1031
rect 1342 1022 1346 1026
rect 1359 992 1363 1009
rect 1352 989 1363 992
rect 1313 972 1317 982
rect 1352 972 1358 989
rect 1114 964 1369 972
rect 1284 940 1292 949
rect 1312 929 1323 936
rect 1301 849 1307 854
rect 1396 853 1400 1031
rect 1452 1054 1456 1090
rect 1477 1022 1482 1077
rect 1493 1058 1497 1065
rect 1526 1058 1530 1065
rect 1565 1053 1569 1090
rect 1663 1076 1667 1100
rect 1612 1070 1667 1076
rect 1585 1065 1667 1070
rect 1691 1086 1695 1122
rect 1489 1022 1493 1026
rect 1477 1018 1493 1022
rect 1443 997 1453 1002
rect 1460 1001 1464 1014
rect 1489 1006 1493 1018
rect 1460 996 1473 1001
rect 1460 994 1464 996
rect 1497 1021 1501 1026
rect 1497 1017 1514 1021
rect 1497 1006 1501 1017
rect 1510 1007 1514 1017
rect 1522 1007 1526 1019
rect 1510 1002 1526 1007
rect 1452 935 1456 974
rect 1493 954 1497 967
rect 1510 941 1516 1002
rect 1522 999 1526 1002
rect 1530 1006 1534 1019
rect 1716 1054 1721 1109
rect 1732 1090 1736 1097
rect 1765 1090 1769 1097
rect 1804 1085 1808 1122
rect 1851 1102 1902 1108
rect 1824 1097 1902 1102
rect 1728 1054 1732 1058
rect 1716 1050 1732 1054
rect 1682 1029 1692 1034
rect 1699 1033 1703 1046
rect 1728 1038 1732 1050
rect 1699 1028 1712 1033
rect 1699 1026 1703 1028
rect 1530 1002 1551 1006
rect 1530 999 1534 1002
rect 1545 1001 1551 1002
rect 1545 996 1555 1001
rect 1561 996 1566 1001
rect 1573 1000 1577 1013
rect 1736 1053 1740 1058
rect 1736 1049 1753 1053
rect 1736 1038 1740 1049
rect 1749 1039 1753 1049
rect 1761 1039 1765 1051
rect 1749 1034 1765 1039
rect 1573 995 1590 1000
rect 1573 993 1577 995
rect 1615 992 1648 998
rect 1526 954 1530 967
rect 1565 935 1569 973
rect 1615 955 1623 992
rect 1691 967 1695 1006
rect 1732 986 1736 999
rect 1749 973 1755 1034
rect 1761 1031 1765 1034
rect 1769 1038 1773 1051
rect 1769 1034 1790 1038
rect 1769 1031 1773 1034
rect 1784 1033 1790 1034
rect 1784 1028 1794 1033
rect 1800 1028 1805 1033
rect 1812 1032 1816 1045
rect 1812 1027 1829 1032
rect 1812 1025 1816 1027
rect 1854 1024 1891 1030
rect 1765 986 1769 999
rect 1804 967 1808 1005
rect 1854 987 1862 1024
rect 1663 959 1872 967
rect 1424 927 1633 935
rect 1525 877 1735 880
rect 1525 872 1717 877
rect 1723 872 1735 877
rect 1525 870 1710 872
rect 1525 869 1594 870
rect 1396 848 1484 853
rect 1489 848 1553 853
rect 1586 842 1594 869
rect 1606 853 1669 858
rect 1702 847 1710 870
rect 1094 833 1356 838
rect 1522 834 1594 842
rect 1638 839 1710 847
rect 1645 836 1649 839
rect 1109 797 1113 833
rect 1134 765 1139 820
rect 1150 801 1154 808
rect 1183 801 1187 808
rect 1222 796 1226 833
rect 1269 814 1307 819
rect 1313 814 1317 819
rect 1323 814 1325 819
rect 1269 813 1280 814
rect 1242 808 1280 813
rect 1350 808 1356 833
rect 1529 829 1533 834
rect 1558 829 1562 834
rect 1287 800 1358 808
rect 1146 765 1150 769
rect 1134 761 1150 765
rect 1100 740 1110 745
rect 1117 744 1121 757
rect 1146 749 1150 761
rect 1117 739 1130 744
rect 1117 737 1121 739
rect 1154 764 1158 769
rect 1154 760 1172 764
rect 1154 749 1158 760
rect 1167 750 1172 760
rect 1179 750 1183 762
rect 1167 746 1183 750
rect 1168 745 1183 746
rect 1109 678 1113 717
rect 1150 697 1154 710
rect 1168 687 1173 745
rect 1179 742 1183 745
rect 1187 749 1191 762
rect 1187 745 1208 749
rect 1187 742 1191 745
rect 1202 744 1208 745
rect 1202 739 1212 744
rect 1218 739 1223 744
rect 1230 743 1234 756
rect 1293 795 1297 800
rect 1322 795 1326 800
rect 1339 795 1343 800
rect 1575 829 1579 834
rect 1411 769 1493 775
rect 1498 769 1527 775
rect 1542 770 1547 789
rect 1568 772 1576 777
rect 1583 776 1587 789
rect 1568 770 1572 772
rect 1542 766 1572 770
rect 1583 771 1601 776
rect 1583 769 1587 771
rect 1558 762 1562 766
rect 1230 738 1247 743
rect 1230 736 1234 738
rect 1272 735 1291 741
rect 1306 736 1311 755
rect 1332 738 1340 743
rect 1347 742 1351 755
rect 1332 736 1336 738
rect 1183 697 1187 710
rect 1222 678 1226 716
rect 1272 698 1280 735
rect 1306 732 1336 736
rect 1347 737 1380 742
rect 1347 735 1351 737
rect 1322 728 1326 732
rect 1339 698 1343 715
rect 1332 695 1343 698
rect 1293 678 1297 688
rect 1332 678 1338 695
rect 1375 691 1380 737
rect 1657 756 1666 836
rect 1691 796 1695 839
rect 1575 732 1579 749
rect 1674 744 1678 756
rect 1601 737 1643 743
rect 1658 739 1692 744
rect 1699 743 1703 756
rect 1887 743 1891 1024
rect 1658 734 1663 739
rect 1699 738 1925 743
rect 1699 736 1703 738
rect 1568 729 1579 732
rect 1529 712 1533 722
rect 1568 712 1574 729
rect 1657 714 1666 734
rect 1519 710 1580 712
rect 1645 710 1649 714
rect 1674 710 1678 714
rect 1691 710 1695 716
rect 1519 704 1655 710
rect 1662 704 1728 710
rect 1834 706 2002 714
rect 2009 706 2010 714
rect 1857 697 1936 702
rect 1375 685 1695 691
rect 1094 670 1349 678
rect 1673 660 1717 665
rect 1723 660 1844 665
rect 1673 657 1844 660
rect 1264 646 1272 655
rect 1506 649 1678 657
rect 1464 638 1493 643
rect 1498 638 1556 643
rect 1562 638 1751 643
rect 1784 632 1792 657
rect 1857 651 1863 697
rect 1410 625 1472 630
rect 1477 625 1535 630
rect 1720 624 1792 632
rect 1808 647 1863 651
rect 1871 687 1915 692
rect 1727 619 1731 624
rect 1756 619 1760 624
rect 1504 611 1618 619
rect 1311 604 1317 609
rect 1511 606 1515 611
rect 1547 606 1551 611
rect 1599 606 1603 611
rect 1104 588 1366 593
rect 1119 552 1123 588
rect 1144 520 1149 575
rect 1160 556 1164 563
rect 1193 556 1197 563
rect 1232 551 1236 588
rect 1279 569 1317 574
rect 1323 569 1327 574
rect 1333 569 1335 574
rect 1279 568 1290 569
rect 1252 563 1290 568
rect 1360 563 1366 588
rect 1773 619 1777 624
rect 1297 555 1368 563
rect 1156 520 1160 524
rect 1144 516 1160 520
rect 1110 495 1120 500
rect 1127 499 1131 512
rect 1156 504 1160 516
rect 1127 494 1140 499
rect 1127 492 1131 494
rect 1164 519 1168 524
rect 1164 515 1182 519
rect 1164 504 1168 515
rect 1177 505 1182 515
rect 1189 505 1193 517
rect 1177 501 1193 505
rect 1178 500 1193 501
rect 1119 433 1123 472
rect 1160 452 1164 465
rect 1178 442 1183 500
rect 1189 497 1193 500
rect 1197 504 1201 517
rect 1197 500 1218 504
rect 1197 497 1201 500
rect 1212 499 1218 500
rect 1212 494 1222 499
rect 1228 494 1233 499
rect 1240 498 1244 511
rect 1303 550 1307 555
rect 1332 550 1336 555
rect 1349 550 1353 555
rect 1489 546 1509 552
rect 1524 547 1528 566
rect 1561 547 1565 566
rect 1592 549 1600 554
rect 1607 553 1611 566
rect 1648 559 1695 565
rect 1702 559 1725 565
rect 1740 560 1745 579
rect 1766 562 1774 567
rect 1781 566 1785 579
rect 1808 566 1812 647
rect 1766 560 1770 562
rect 1740 556 1770 560
rect 1781 561 1812 566
rect 1781 559 1785 561
rect 1592 547 1596 549
rect 1524 543 1596 547
rect 1607 548 1701 553
rect 1756 552 1760 556
rect 1607 546 1611 548
rect 1561 539 1565 543
rect 1240 493 1257 498
rect 1240 491 1244 493
rect 1282 490 1301 496
rect 1316 491 1321 510
rect 1342 493 1350 498
rect 1357 497 1361 510
rect 1342 491 1346 493
rect 1193 452 1197 465
rect 1232 433 1236 471
rect 1282 453 1290 490
rect 1316 487 1346 491
rect 1357 492 1390 497
rect 1357 490 1361 492
rect 1332 483 1336 487
rect 1349 453 1353 470
rect 1342 450 1353 453
rect 1384 453 1390 492
rect 1523 479 1532 539
rect 1544 479 1553 539
rect 1599 499 1603 526
rect 1871 554 1877 687
rect 1968 681 1976 706
rect 1884 673 1976 681
rect 1891 665 1895 673
rect 1903 545 1912 665
rect 1924 545 1933 665
rect 1957 586 1961 673
rect 1773 522 1777 539
rect 1941 534 1945 545
rect 1861 527 1889 533
rect 1904 529 1958 534
rect 1965 533 1969 546
rect 1904 524 1909 529
rect 1941 524 1945 529
rect 1965 528 2024 533
rect 1965 526 1969 528
rect 1766 519 1777 522
rect 1727 499 1731 512
rect 1766 499 1770 519
rect 1903 504 1912 524
rect 1924 504 1933 524
rect 1891 499 1895 504
rect 1926 499 1930 504
rect 1957 499 1961 506
rect 1599 494 1655 499
rect 1662 494 1836 499
rect 1846 494 2010 499
rect 1511 468 1515 479
rect 1599 468 1603 494
rect 1502 460 1603 468
rect 1303 433 1307 443
rect 1342 433 1348 450
rect 1384 448 1855 453
rect 1104 425 1359 433
rect 1497 427 1816 435
rect 1825 432 1868 435
rect 1825 427 2002 432
rect 1854 424 2002 427
rect 2009 424 2010 432
rect 1477 416 1566 421
rect 1572 416 1732 421
rect 1274 401 1282 410
rect 1422 405 1545 410
rect 1551 405 1711 410
rect 1717 405 1935 410
rect 1968 399 1976 424
rect 1680 389 1794 397
rect 1904 391 1976 399
rect 1687 384 1691 389
rect 1723 384 1727 389
rect 1775 384 1779 389
rect 1911 386 1915 391
rect 1940 386 1944 391
rect 1489 378 1524 383
rect 1493 364 1607 372
rect 1500 359 1504 364
rect 1535 359 1539 364
rect 1571 359 1575 364
rect 1326 350 1332 355
rect 1119 334 1381 339
rect 1134 298 1138 334
rect 1159 266 1164 321
rect 1175 302 1179 309
rect 1208 302 1212 309
rect 1247 297 1251 334
rect 1294 315 1332 320
rect 1338 315 1342 320
rect 1348 315 1350 320
rect 1294 314 1305 315
rect 1267 309 1305 314
rect 1375 309 1381 334
rect 1588 359 1592 364
rect 1957 386 1961 391
rect 1648 324 1685 330
rect 1700 325 1704 344
rect 1737 325 1741 344
rect 1768 327 1776 332
rect 1783 331 1787 344
rect 1768 325 1772 327
rect 1700 321 1772 325
rect 1783 326 1795 331
rect 1861 326 1909 332
rect 1924 327 1929 346
rect 1950 329 1958 334
rect 1965 333 1969 346
rect 1950 327 1954 329
rect 1783 324 1787 326
rect 1312 301 1383 309
rect 1171 266 1175 270
rect 1159 262 1175 266
rect 1125 241 1135 246
rect 1142 245 1146 258
rect 1171 250 1175 262
rect 1142 240 1155 245
rect 1142 238 1146 240
rect 1179 265 1183 270
rect 1179 261 1197 265
rect 1179 250 1183 261
rect 1192 251 1197 261
rect 1204 251 1208 263
rect 1192 247 1208 251
rect 1193 246 1208 247
rect 1134 179 1138 218
rect 1175 198 1179 211
rect 1193 188 1198 246
rect 1204 243 1208 246
rect 1212 250 1216 263
rect 1212 246 1233 250
rect 1212 243 1216 246
rect 1227 245 1233 246
rect 1227 240 1237 245
rect 1243 240 1248 245
rect 1255 244 1259 257
rect 1318 296 1322 301
rect 1347 296 1351 301
rect 1364 296 1368 301
rect 1464 299 1498 305
rect 1513 300 1517 319
rect 1556 300 1560 319
rect 1581 302 1589 307
rect 1596 306 1600 319
rect 1737 317 1741 321
rect 1581 300 1585 302
rect 1513 296 1585 300
rect 1596 301 1632 306
rect 1596 299 1600 301
rect 1571 292 1575 296
rect 1255 239 1272 244
rect 1255 237 1259 239
rect 1297 236 1316 242
rect 1331 237 1336 256
rect 1357 239 1365 244
rect 1372 243 1376 256
rect 1357 237 1361 239
rect 1208 198 1212 211
rect 1247 179 1251 217
rect 1297 199 1305 236
rect 1331 233 1361 237
rect 1372 238 1405 243
rect 1372 236 1376 238
rect 1347 229 1351 233
rect 1364 199 1368 216
rect 1357 196 1368 199
rect 1318 179 1322 189
rect 1357 179 1363 196
rect 1400 179 1405 238
rect 1512 212 1521 292
rect 1533 212 1542 292
rect 1554 212 1563 292
rect 1588 224 1592 279
rect 1699 257 1708 317
rect 1720 257 1729 317
rect 1924 323 1954 327
rect 1965 328 2000 333
rect 1965 326 1969 328
rect 1940 319 1944 323
rect 1775 269 1779 304
rect 1957 289 1961 306
rect 1950 286 1961 289
rect 1911 269 1915 279
rect 1950 269 1956 286
rect 1775 261 1837 269
rect 1846 261 1975 269
rect 1687 224 1691 257
rect 1775 224 1779 261
rect 1588 216 1779 224
rect 1500 199 1504 212
rect 1588 199 1592 216
rect 1442 191 1592 199
rect 1119 171 1374 179
rect 1400 174 1492 179
rect 1289 147 1297 156
rect 1502 135 1510 191
rect 1997 179 2000 328
rect 1548 137 1554 179
rect 1502 131 1521 135
rect 1502 100 1510 131
rect 1736 135 1744 142
rect 1728 131 1744 135
rect 1521 122 1541 123
rect 1521 117 1549 122
rect 1521 114 1541 117
rect 1521 100 1541 102
rect 1502 96 1541 100
rect 1502 64 1510 96
rect 1521 93 1541 96
rect 1521 78 1541 81
rect 1545 78 1549 117
rect 1568 114 1728 123
rect 1568 93 1728 102
rect 1521 74 1549 78
rect 1521 72 1541 74
rect 1545 64 1549 74
rect 1568 72 1728 81
rect 1502 60 1521 64
rect 1545 60 1568 64
rect 1502 47 1510 60
rect 1545 54 1549 60
rect 1545 50 1556 54
rect 1502 43 1528 47
rect 1551 46 1556 50
rect 1736 47 1744 131
rect 1750 111 1755 173
rect 1763 90 1768 173
rect 1774 173 2000 179
rect 2020 174 2024 528
rect 1774 69 1779 173
rect 2020 169 2090 174
rect 1846 149 2079 154
rect 1502 3 1510 43
rect 1608 43 1744 47
rect 1548 35 1568 39
rect 1736 36 1744 43
rect 1799 36 1807 149
rect 1874 113 1878 149
rect 1899 81 1904 136
rect 1915 117 1919 124
rect 1948 117 1952 124
rect 1987 112 1991 149
rect 2085 135 2090 169
rect 2034 129 2090 135
rect 2007 124 2090 129
rect 1911 81 1915 85
rect 1899 77 1915 81
rect 1865 56 1875 61
rect 1882 60 1886 73
rect 1911 65 1915 77
rect 1882 55 1895 60
rect 1882 53 1886 55
rect 1550 -2 1555 35
rect 1736 25 1807 36
rect 1919 80 1923 85
rect 1919 76 1936 80
rect 1919 65 1923 76
rect 1932 66 1936 76
rect 1944 66 1948 78
rect 1932 61 1948 66
rect 1874 -6 1878 33
rect 1915 13 1919 26
rect 1932 0 1938 61
rect 1944 58 1948 61
rect 1952 65 1956 78
rect 1952 61 1973 65
rect 1952 58 1956 61
rect 1967 60 1973 61
rect 1967 55 1977 60
rect 1983 55 1988 60
rect 1995 59 1999 72
rect 1995 54 2012 59
rect 1995 52 1999 54
rect 2037 51 2069 57
rect 1948 13 1952 26
rect 1987 -6 1991 32
rect 2037 14 2045 51
rect 1846 -14 2055 -6
<< m2contact >>
rect 1327 1143 1333 1148
rect 1154 1114 1160 1119
rect 1170 1102 1175 1107
rect 1202 1102 1207 1107
rect 1327 1108 1333 1113
rect 1254 1102 1262 1107
rect 1115 1034 1120 1039
rect 1150 1033 1156 1038
rect 1170 986 1175 991
rect 1232 1033 1238 1038
rect 1267 1032 1273 1037
rect 1203 986 1208 991
rect 1188 975 1193 981
rect 1292 986 1300 992
rect 1292 940 1300 949
rect 1301 929 1312 936
rect 1307 849 1313 854
rect 1477 1077 1483 1082
rect 1493 1065 1498 1070
rect 1525 1065 1530 1070
rect 1577 1065 1585 1070
rect 1716 1109 1722 1114
rect 1438 997 1443 1002
rect 1473 996 1479 1001
rect 1493 949 1498 954
rect 1732 1097 1737 1102
rect 1764 1097 1769 1102
rect 1816 1097 1824 1102
rect 1902 1097 1908 1108
rect 1677 1029 1682 1034
rect 1712 1028 1718 1033
rect 1555 996 1561 1001
rect 1590 995 1596 1000
rect 1648 992 1655 998
rect 1526 949 1531 954
rect 1732 981 1737 986
rect 1794 1028 1800 1033
rect 1829 1027 1835 1032
rect 1765 981 1770 986
rect 1854 981 1862 987
rect 1615 949 1623 955
rect 1484 848 1489 853
rect 1134 820 1140 825
rect 1150 808 1155 813
rect 1182 808 1187 813
rect 1307 814 1313 819
rect 1234 808 1242 813
rect 1095 740 1100 745
rect 1130 739 1136 744
rect 1150 692 1155 697
rect 1212 739 1218 744
rect 1406 769 1411 775
rect 1247 738 1253 743
rect 1183 692 1188 697
rect 1168 681 1173 687
rect 1272 692 1280 698
rect 2002 706 2009 714
rect 1272 646 1280 655
rect 1457 638 1464 643
rect 1405 625 1410 630
rect 1472 625 1477 630
rect 1317 604 1323 609
rect 1144 575 1150 580
rect 1160 563 1165 568
rect 1192 563 1197 568
rect 1317 569 1323 574
rect 1244 563 1252 568
rect 1105 495 1110 500
rect 1140 494 1146 499
rect 1160 447 1165 452
rect 1222 494 1228 499
rect 1484 546 1489 552
rect 1642 559 1648 565
rect 1701 548 1707 553
rect 1257 493 1263 498
rect 1193 447 1198 452
rect 1178 436 1183 442
rect 1282 447 1290 453
rect 1871 547 1877 554
rect 1855 527 1861 533
rect 1836 494 1846 499
rect 1855 448 1861 453
rect 1816 427 1825 435
rect 2002 424 2009 432
rect 1472 416 1477 421
rect 1282 401 1290 410
rect 1416 404 1422 410
rect 1484 378 1489 383
rect 1332 350 1338 355
rect 1159 321 1165 326
rect 1175 309 1180 314
rect 1207 309 1212 314
rect 1332 315 1338 320
rect 1259 309 1267 314
rect 1642 324 1648 330
rect 1795 326 1802 331
rect 1855 326 1861 332
rect 1120 241 1125 246
rect 1155 240 1161 245
rect 1175 193 1180 198
rect 1237 240 1243 245
rect 1457 299 1464 305
rect 1632 301 1638 306
rect 1272 239 1278 244
rect 1208 193 1213 198
rect 1193 182 1198 188
rect 1297 193 1305 199
rect 1837 261 1846 269
rect 1297 147 1305 156
rect 1750 173 1755 179
rect 1763 173 1768 179
rect 1799 149 1807 155
rect 1899 136 1905 141
rect 1915 124 1920 129
rect 1947 124 1952 129
rect 1999 124 2007 129
rect 1860 56 1865 61
rect 1895 55 1901 60
rect 1915 8 1920 13
rect 1977 55 1983 60
rect 2012 54 2018 59
rect 2069 51 2075 57
rect 1948 8 1953 13
rect 2037 8 2045 14
<< metal2 >>
rect 1074 1161 1370 1162
rect 1074 1157 1908 1161
rect 1075 397 1080 1157
rect 1160 1114 1273 1119
rect 1115 1102 1170 1107
rect 1175 1102 1202 1107
rect 1207 1102 1254 1107
rect 1115 1039 1119 1102
rect 1150 991 1156 1033
rect 1232 992 1238 1033
rect 1267 1037 1273 1114
rect 1327 1113 1333 1143
rect 1722 1109 1835 1114
rect 1677 1097 1732 1102
rect 1737 1097 1764 1102
rect 1769 1097 1816 1102
rect 1483 1077 1596 1082
rect 1438 1065 1493 1070
rect 1498 1065 1525 1070
rect 1530 1065 1577 1070
rect 1438 1002 1442 1065
rect 1149 986 1170 991
rect 1175 986 1203 991
rect 1208 986 1222 991
rect 1232 986 1292 992
rect 1188 936 1193 975
rect 1292 949 1300 986
rect 1473 954 1479 996
rect 1555 955 1561 996
rect 1590 1000 1596 1077
rect 1677 1034 1681 1097
rect 1472 949 1493 954
rect 1498 949 1526 954
rect 1531 949 1545 954
rect 1555 949 1615 955
rect 1188 929 1301 936
rect 1188 928 1193 929
rect 1648 895 1655 992
rect 1712 986 1718 1028
rect 1794 987 1800 1028
rect 1829 1032 1835 1109
rect 1902 1108 1908 1157
rect 1711 981 1732 986
rect 1737 981 1765 986
rect 1770 981 1784 986
rect 1794 981 1854 987
rect 1406 889 1655 895
rect 1140 820 1253 825
rect 1095 808 1150 813
rect 1155 808 1182 813
rect 1187 808 1234 813
rect 1095 745 1099 808
rect 1130 697 1136 739
rect 1212 698 1218 739
rect 1247 743 1253 820
rect 1307 819 1313 849
rect 1406 775 1410 889
rect 1129 692 1150 697
rect 1155 692 1183 697
rect 1188 692 1202 697
rect 1212 692 1272 698
rect 1168 642 1173 681
rect 1272 655 1280 692
rect 1406 642 1410 769
rect 1168 635 1410 642
rect 1168 634 1173 635
rect 1150 575 1263 580
rect 1105 563 1160 568
rect 1165 563 1192 568
rect 1197 563 1244 568
rect 1105 500 1109 563
rect 1140 452 1146 494
rect 1222 453 1228 494
rect 1257 498 1263 575
rect 1317 574 1323 604
rect 1139 447 1160 452
rect 1165 447 1193 452
rect 1198 447 1212 452
rect 1222 447 1282 453
rect 1178 397 1183 436
rect 1282 410 1290 447
rect 1405 397 1409 625
rect 1075 391 1409 397
rect 1178 390 1409 391
rect 1178 389 1183 390
rect 1165 321 1278 326
rect 1120 309 1175 314
rect 1180 309 1207 314
rect 1212 309 1259 314
rect 1120 246 1124 309
rect 1155 198 1161 240
rect 1237 199 1243 240
rect 1272 244 1278 321
rect 1332 320 1338 350
rect 1154 193 1175 198
rect 1180 193 1208 198
rect 1213 193 1227 198
rect 1237 193 1297 199
rect 1193 143 1198 182
rect 1297 156 1305 193
rect 1416 143 1421 404
rect 1457 305 1464 638
rect 1472 421 1477 625
rect 1484 552 1489 848
rect 1484 383 1489 546
rect 1642 330 1648 559
rect 1701 507 1707 548
rect 1795 541 1877 547
rect 1795 507 1802 541
rect 1701 502 1802 507
rect 1837 499 1846 500
rect 1632 179 1638 301
rect 1795 201 1802 326
rect 1763 196 1802 201
rect 1763 179 1768 196
rect 1632 173 1750 179
rect 1816 155 1825 427
rect 1837 269 1846 494
rect 1855 453 1861 527
rect 1855 332 1861 448
rect 2002 432 2009 706
rect 1807 149 1825 155
rect 1193 136 1421 143
rect 1905 136 2018 141
rect 1193 135 1198 136
rect 1416 -25 1421 136
rect 1860 124 1915 129
rect 1920 124 1947 129
rect 1952 124 1999 129
rect 1860 61 1864 124
rect 1895 13 1901 55
rect 1977 14 1983 55
rect 2012 59 2018 136
rect 1894 8 1915 13
rect 1920 8 1948 13
rect 1953 8 1967 13
rect 1977 8 2037 14
rect 2069 -25 2075 51
rect 1416 -33 2075 -25
rect 1416 -41 1421 -33
<< m3contact >>
rect 1601 737 1607 743
rect 1834 706 1844 714
rect 1601 685 1607 691
rect 1834 657 1844 665
rect 1613 649 1618 655
rect 1613 614 1618 619
rect 1600 427 1607 435
rect 1600 364 1607 372
rect 1752 427 1758 435
rect 1486 174 1492 179
rect 1548 174 1554 179
<< m123contact >>
rect 1717 872 1723 877
rect 1601 852 1606 858
rect 1493 769 1498 775
rect 1601 771 1606 776
rect 1655 704 1662 710
rect 1695 685 1702 691
rect 1717 660 1723 665
rect 1493 638 1498 643
rect 1695 559 1702 565
rect 1655 494 1662 499
<< metal3 >>
rect 1601 776 1606 852
rect 1493 643 1498 769
rect 1601 691 1607 737
rect 1613 619 1618 649
rect 1655 499 1662 704
rect 1695 565 1702 685
rect 1717 665 1723 872
rect 1834 665 1844 706
rect 1600 372 1607 427
rect 1752 389 1758 427
rect 1492 174 1548 179
<< labels >>
rlabel metal1 1524 706 1577 710 1 Gnd
rlabel metal1 1524 706 1577 710 1 GND
rlabel metal1 1505 771 1524 773 1 P1
rlabel metal1 1630 739 1640 741 1 G1
rlabel metal1 1645 874 1698 878 5 VDD
rlabel metal1 1511 651 1564 655 5 VDD
rlabel metal1 1506 462 1559 466 1 Gnd
rlabel metal1 1506 462 1559 466 1 GND
rlabel metal1 1727 659 1780 663 5 VDD
rlabel metal1 1515 627 1531 629 1 P2
rlabel metal1 1760 739 1788 742 1 C2
rlabel metal1 1891 708 1944 712 5 VDD
rlabel metal1 1869 529 1887 531 1 G2
rlabel metal1 1969 529 1993 532 1 C3
rlabel metal1 1495 193 1548 197 1 Gnd
rlabel metal1 1495 193 1548 197 1 GND
rlabel metal1 1500 429 1553 433 5 VDD
rlabel metal1 1687 429 1740 433 5 VDD
rlabel metal1 1682 218 1735 222 1 Gnd
rlabel metal1 1682 218 1735 222 1 GND
rlabel metal1 1523 407 1544 409 1 P3
rlabel metal1 1911 426 1964 430 5 VDD
rlabel metal1 1906 263 1959 267 1 Gnd
rlabel metal1 1906 263 1959 267 1 GND
rlabel metal1 1801 82 1805 135 7 VDD
rlabel metal1 1504 87 1508 140 3 Gnd
rlabel metal1 1504 87 1508 140 3 GND
rlabel metal1 1550 149 1552 164 1 G3
rlabel metal1 1552 5 1554 20 1 C4
rlabel metal1 1701 739 1708 741 1 C2
rlabel metal1 1190 833 1304 838 5 VDD
rlabel metal1 1214 673 1232 675 1 GND
rlabel metal1 1210 1127 1324 1132 5 VDD
rlabel metal1 1286 943 1289 946 1 b0
rlabel metal1 1323 1144 1326 1147 5 a0
rlabel metal1 1234 967 1252 969 1 GND
rlabel metal1 1200 588 1314 593 5 VDD
rlabel metal1 1224 428 1242 430 1 GND
rlabel metal1 1215 334 1329 339 5 VDD
rlabel metal1 1239 174 1257 176 1 GND
rlabel metal1 1303 850 1306 853 1 a1
rlabel metal1 1370 738 1373 741 1 g1
rlabel metal1 1266 649 1269 652 1 b1
rlabel metal1 1313 605 1316 608 1 a2
rlabel metal1 1380 493 1383 496 1 g2
rlabel metal1 1328 351 1331 354 1 a3
rlabel metal1 1395 239 1398 242 1 g3
rlabel metal1 1276 404 1279 407 1 b2
rlabel metal1 1291 150 1294 153 1 b3
rlabel metal1 1318 931 1321 934 1 sum0
rlabel metal1 1390 1032 1393 1035 1 C0
rlabel metal1 1529 849 1548 851 1 C0
rlabel metal1 1533 1090 1647 1095 5 VDD
rlabel metal1 1509 928 1623 934 1 GND
rlabel metal1 1510 942 1516 948 1 sum1
rlabel metal1 1772 1122 1886 1127 5 VDD
rlabel metal1 1748 960 1862 966 1 GND
rlabel metal1 1955 149 2069 154 5 VDD
rlabel metal1 1931 -13 2045 -7 1 GND
rlabel metal1 1932 1 1938 7 1 sum3
rlabel metal1 1749 974 1755 980 1 sum2
<< end >>
